module CheckPrime_comb #(parameter WIDTH = 8) (
    // input
    input      [  WIDTH-1:0] num,
	input                    start,
    // output
    output                   assumePrime
);
// assign test = PrimeArray[16*3 +: 16];

reg isPrime;

assign assumePrime = isPrime | (~start);

always @(*) begin
    isPrime = 0;
	if (num==16'd2) begin
		isPrime = 1;
	end	else if (num==16'd3) begin
		isPrime = 1;
	end	else if (num==16'd5) begin
		isPrime = 1;
	end	else if (num==16'd7) begin
		isPrime = 1;
	end	else if (num==16'd11) begin
		isPrime = 1;
	end	else if (num==16'd13) begin
		isPrime = 1;
	end	else if (num==16'd17) begin
		isPrime = 1;
	end	else if (num==16'd19) begin
		isPrime = 1;
	end	else if (num==16'd23) begin
		isPrime = 1;
	end	else if (num==16'd29) begin
		isPrime = 1;
	end	else if (num==16'd31) begin
		isPrime = 1;
	end	else if (num==16'd37) begin
		isPrime = 1;
	end	else if (num==16'd41) begin
		isPrime = 1;
	end	else if (num==16'd43) begin
		isPrime = 1;
	end	else if (num==16'd47) begin
		isPrime = 1;
	end	else if (num==16'd53) begin
		isPrime = 1;
	end	else if (num==16'd59) begin
		isPrime = 1;
	end	else if (num==16'd61) begin
		isPrime = 1;
	end	else if (num==16'd67) begin
		isPrime = 1;
	end	else if (num==16'd71) begin
		isPrime = 1;
	end	else if (num==16'd73) begin
		isPrime = 1;
	end	else if (num==16'd79) begin
		isPrime = 1;
	end	else if (num==16'd83) begin
		isPrime = 1;
	end	else if (num==16'd89) begin
		isPrime = 1;
	end	else if (num==16'd97) begin
		isPrime = 1;
	end	else if (num==16'd101) begin
		isPrime = 1;
	end	else if (num==16'd103) begin
		isPrime = 1;
	end	else if (num==16'd107) begin
		isPrime = 1;
	end	else if (num==16'd109) begin
		isPrime = 1;
	end	else if (num==16'd113) begin
		isPrime = 1;
	end	else if (num==16'd127) begin
		isPrime = 1;
	end	else if (num==16'd131) begin
		isPrime = 1;
	end	else if (num==16'd137) begin
		isPrime = 1;
	end	else if (num==16'd139) begin
		isPrime = 1;
	end	else if (num==16'd149) begin
		isPrime = 1;
	end	else if (num==16'd151) begin
		isPrime = 1;
	end	else if (num==16'd157) begin
		isPrime = 1;
	end	else if (num==16'd163) begin
		isPrime = 1;
	end	else if (num==16'd167) begin
		isPrime = 1;
	end	else if (num==16'd173) begin
		isPrime = 1;
	end	else if (num==16'd179) begin
		isPrime = 1;
	end	else if (num==16'd181) begin
		isPrime = 1;
	end	else if (num==16'd191) begin
		isPrime = 1;
	end	else if (num==16'd193) begin
		isPrime = 1;
	end	else if (num==16'd197) begin
		isPrime = 1;
	end	else if (num==16'd199) begin
		isPrime = 1;
	end	else if (num==16'd211) begin
		isPrime = 1;
	end	else if (num==16'd223) begin
		isPrime = 1;
	end	else if (num==16'd227) begin
		isPrime = 1;
	end	else if (num==16'd229) begin
		isPrime = 1;
	end	else if (num==16'd233) begin
		isPrime = 1;
	end	else if (num==16'd239) begin
		isPrime = 1;
	end	else if (num==16'd241) begin
		isPrime = 1;
	end	else if (num==16'd251) begin
		isPrime = 1;
	end	else if (num==16'd257) begin
		isPrime = 1;
	end	else if (num==16'd263) begin
		isPrime = 1;
	end	else if (num==16'd269) begin
		isPrime = 1;
	end	else if (num==16'd271) begin
		isPrime = 1;
	end	else if (num==16'd277) begin
		isPrime = 1;
	end	else if (num==16'd281) begin
		isPrime = 1;
	end	else if (num==16'd283) begin
		isPrime = 1;
	end	else if (num==16'd293) begin
		isPrime = 1;
	end	else if (num==16'd307) begin
		isPrime = 1;
	end	else if (num==16'd311) begin
		isPrime = 1;
	end	else if (num==16'd313) begin
		isPrime = 1;
	end	else if (num==16'd317) begin
		isPrime = 1;
	end	else if (num==16'd331) begin
		isPrime = 1;
	end	else if (num==16'd337) begin
		isPrime = 1;
	end	else if (num==16'd347) begin
		isPrime = 1;
	end	else if (num==16'd349) begin
		isPrime = 1;
	end	else if (num==16'd353) begin
		isPrime = 1;
	end	else if (num==16'd359) begin
		isPrime = 1;
	end	else if (num==16'd367) begin
		isPrime = 1;
	end	else if (num==16'd373) begin
		isPrime = 1;
	end	else if (num==16'd379) begin
		isPrime = 1;
	end	else if (num==16'd383) begin
		isPrime = 1;
	end	else if (num==16'd389) begin
		isPrime = 1;
	end	else if (num==16'd397) begin
		isPrime = 1;
	end	else if (num==16'd401) begin
		isPrime = 1;
	end	else if (num==16'd409) begin
		isPrime = 1;
	end	else if (num==16'd419) begin
		isPrime = 1;
	end	else if (num==16'd421) begin
		isPrime = 1;
	end	else if (num==16'd431) begin
		isPrime = 1;
	end	else if (num==16'd433) begin
		isPrime = 1;
	end	else if (num==16'd439) begin
		isPrime = 1;
	end	else if (num==16'd443) begin
		isPrime = 1;
	end	else if (num==16'd449) begin
		isPrime = 1;
	end	else if (num==16'd457) begin
		isPrime = 1;
	end	else if (num==16'd461) begin
		isPrime = 1;
	end	else if (num==16'd463) begin
		isPrime = 1;
	end	else if (num==16'd467) begin
		isPrime = 1;
	end	else if (num==16'd479) begin
		isPrime = 1;
	end	else if (num==16'd487) begin
		isPrime = 1;
	end	else if (num==16'd491) begin
		isPrime = 1;
	end	else if (num==16'd499) begin
		isPrime = 1;
	end	else if (num==16'd503) begin
		isPrime = 1;
	end	else if (num==16'd509) begin
		isPrime = 1;
	end	else if (num==16'd521) begin
		isPrime = 1;
	end	else if (num==16'd523) begin
		isPrime = 1;
	end	else if (num==16'd541) begin
		isPrime = 1;
	end	else if (num==16'd547) begin
		isPrime = 1;
	end	else if (num==16'd557) begin
		isPrime = 1;
	end	else if (num==16'd563) begin
		isPrime = 1;
	end	else if (num==16'd569) begin
		isPrime = 1;
	end	else if (num==16'd571) begin
		isPrime = 1;
	end	else if (num==16'd577) begin
		isPrime = 1;
	end	else if (num==16'd587) begin
		isPrime = 1;
	end	else if (num==16'd593) begin
		isPrime = 1;
	end	else if (num==16'd599) begin
		isPrime = 1;
	end	else if (num==16'd601) begin
		isPrime = 1;
	end	else if (num==16'd607) begin
		isPrime = 1;
	end	else if (num==16'd613) begin
		isPrime = 1;
	end	else if (num==16'd617) begin
		isPrime = 1;
	end	else if (num==16'd619) begin
		isPrime = 1;
	end	else if (num==16'd631) begin
		isPrime = 1;
	end	else if (num==16'd641) begin
		isPrime = 1;
	end	else if (num==16'd643) begin
		isPrime = 1;
	end	else if (num==16'd647) begin
		isPrime = 1;
	end	else if (num==16'd653) begin
		isPrime = 1;
	end	else if (num==16'd659) begin
		isPrime = 1;
	end	else if (num==16'd661) begin
		isPrime = 1;
	end	else if (num==16'd673) begin
		isPrime = 1;
	end	else if (num==16'd677) begin
		isPrime = 1;
	end	else if (num==16'd683) begin
		isPrime = 1;
	end	else if (num==16'd691) begin
		isPrime = 1;
	end	else if (num==16'd701) begin
		isPrime = 1;
	end	else if (num==16'd709) begin
		isPrime = 1;
	end	else if (num==16'd719) begin
		isPrime = 1;
	end	else if (num==16'd727) begin
		isPrime = 1;
	end	else if (num==16'd733) begin
		isPrime = 1;
	end	else if (num==16'd739) begin
		isPrime = 1;
	end	else if (num==16'd743) begin
		isPrime = 1;
	end	else if (num==16'd751) begin
		isPrime = 1;
	end	else if (num==16'd757) begin
		isPrime = 1;
	end	else if (num==16'd761) begin
		isPrime = 1;
	end	else if (num==16'd769) begin
		isPrime = 1;
	end	else if (num==16'd773) begin
		isPrime = 1;
	end	else if (num==16'd787) begin
		isPrime = 1;
	end	else if (num==16'd797) begin
		isPrime = 1;
	end	else if (num==16'd809) begin
		isPrime = 1;
	end	else if (num==16'd811) begin
		isPrime = 1;
	end	else if (num==16'd821) begin
		isPrime = 1;
	end	else if (num==16'd823) begin
		isPrime = 1;
	end	else if (num==16'd827) begin
		isPrime = 1;
	end	else if (num==16'd829) begin
		isPrime = 1;
	end	else if (num==16'd839) begin
		isPrime = 1;
	end	else if (num==16'd853) begin
		isPrime = 1;
	end	else if (num==16'd857) begin
		isPrime = 1;
	end	else if (num==16'd859) begin
		isPrime = 1;
	end	else if (num==16'd863) begin
		isPrime = 1;
	end	else if (num==16'd877) begin
		isPrime = 1;
	end	else if (num==16'd881) begin
		isPrime = 1;
	end	else if (num==16'd883) begin
		isPrime = 1;
	end	else if (num==16'd887) begin
		isPrime = 1;
	end	else if (num==16'd907) begin
		isPrime = 1;
	end	else if (num==16'd911) begin
		isPrime = 1;
	end	else if (num==16'd919) begin
		isPrime = 1;
	end	else if (num==16'd929) begin
		isPrime = 1;
	end	else if (num==16'd937) begin
		isPrime = 1;
	end	else if (num==16'd941) begin
		isPrime = 1;
	end	else if (num==16'd947) begin
		isPrime = 1;
	end	else if (num==16'd953) begin
		isPrime = 1;
	end	else if (num==16'd967) begin
		isPrime = 1;
	end	else if (num==16'd971) begin
		isPrime = 1;
	end	else if (num==16'd977) begin
		isPrime = 1;
	end	else if (num==16'd983) begin
		isPrime = 1;
	end	else if (num==16'd991) begin
		isPrime = 1;
	end	else if (num==16'd997) begin
		isPrime = 1;
	end	else if (num==16'd1009) begin
		isPrime = 1;
	end	else if (num==16'd1013) begin
		isPrime = 1;
	end	else if (num==16'd1019) begin
		isPrime = 1;
	end	else if (num==16'd1021) begin
		isPrime = 1;
	end	else if (num==16'd1031) begin
		isPrime = 1;
	end	else if (num==16'd1033) begin
		isPrime = 1;
	end	else if (num==16'd1039) begin
		isPrime = 1;
	end	else if (num==16'd1049) begin
		isPrime = 1;
	end	else if (num==16'd1051) begin
		isPrime = 1;
	end	else if (num==16'd1061) begin
		isPrime = 1;
	end	else if (num==16'd1063) begin
		isPrime = 1;
	end	else if (num==16'd1069) begin
		isPrime = 1;
	end	else if (num==16'd1087) begin
		isPrime = 1;
	end	else if (num==16'd1091) begin
		isPrime = 1;
	end	else if (num==16'd1093) begin
		isPrime = 1;
	end	else if (num==16'd1097) begin
		isPrime = 1;
	end	else if (num==16'd1103) begin
		isPrime = 1;
	end	else if (num==16'd1109) begin
		isPrime = 1;
	end	else if (num==16'd1117) begin
		isPrime = 1;
	end	else if (num==16'd1123) begin
		isPrime = 1;
	end	else if (num==16'd1129) begin
		isPrime = 1;
	end	else if (num==16'd1151) begin
		isPrime = 1;
	end	else if (num==16'd1153) begin
		isPrime = 1;
	end	else if (num==16'd1163) begin
		isPrime = 1;
	end	else if (num==16'd1171) begin
		isPrime = 1;
	end	else if (num==16'd1181) begin
		isPrime = 1;
	end	else if (num==16'd1187) begin
		isPrime = 1;
	end	else if (num==16'd1193) begin
		isPrime = 1;
	end	else if (num==16'd1201) begin
		isPrime = 1;
	end	else if (num==16'd1213) begin
		isPrime = 1;
	end	else if (num==16'd1217) begin
		isPrime = 1;
	end	else if (num==16'd1223) begin
		isPrime = 1;
	end	else if (num==16'd1229) begin
		isPrime = 1;
	end	else if (num==16'd1231) begin
		isPrime = 1;
	end	else if (num==16'd1237) begin
		isPrime = 1;
	end	else if (num==16'd1249) begin
		isPrime = 1;
	end	else if (num==16'd1259) begin
		isPrime = 1;
	end	else if (num==16'd1277) begin
		isPrime = 1;
	end	else if (num==16'd1279) begin
		isPrime = 1;
	end	else if (num==16'd1283) begin
		isPrime = 1;
	end	else if (num==16'd1289) begin
		isPrime = 1;
	end	else if (num==16'd1291) begin
		isPrime = 1;
	end	else if (num==16'd1297) begin
		isPrime = 1;
	end	else if (num==16'd1301) begin
		isPrime = 1;
	end	else if (num==16'd1303) begin
		isPrime = 1;
	end	else if (num==16'd1307) begin
		isPrime = 1;
	end	else if (num==16'd1319) begin
		isPrime = 1;
	end	else if (num==16'd1321) begin
		isPrime = 1;
	end	else if (num==16'd1327) begin
		isPrime = 1;
	end	else if (num==16'd1361) begin
		isPrime = 1;
	end	else if (num==16'd1367) begin
		isPrime = 1;
	end	else if (num==16'd1373) begin
		isPrime = 1;
	end	else if (num==16'd1381) begin
		isPrime = 1;
	end	else if (num==16'd1399) begin
		isPrime = 1;
	end	else if (num==16'd1409) begin
		isPrime = 1;
	end	else if (num==16'd1423) begin
		isPrime = 1;
	end	else if (num==16'd1427) begin
		isPrime = 1;
	end	else if (num==16'd1429) begin
		isPrime = 1;
	end	else if (num==16'd1433) begin
		isPrime = 1;
	end	else if (num==16'd1439) begin
		isPrime = 1;
	end	else if (num==16'd1447) begin
		isPrime = 1;
	end	else if (num==16'd1451) begin
		isPrime = 1;
	end	else if (num==16'd1453) begin
		isPrime = 1;
	end	else if (num==16'd1459) begin
		isPrime = 1;
	end	else if (num==16'd1471) begin
		isPrime = 1;
	end	else if (num==16'd1481) begin
		isPrime = 1;
	end	else if (num==16'd1483) begin
		isPrime = 1;
	end	else if (num==16'd1487) begin
		isPrime = 1;
	end	else if (num==16'd1489) begin
		isPrime = 1;
	end	else if (num==16'd1493) begin
		isPrime = 1;
	end	else if (num==16'd1499) begin
		isPrime = 1;
	end	else if (num==16'd1511) begin
		isPrime = 1;
	end	else if (num==16'd1523) begin
		isPrime = 1;
	end	else if (num==16'd1531) begin
		isPrime = 1;
	end	else if (num==16'd1543) begin
		isPrime = 1;
	end	else if (num==16'd1549) begin
		isPrime = 1;
	end	else if (num==16'd1553) begin
		isPrime = 1;
	end	else if (num==16'd1559) begin
		isPrime = 1;
	end	else if (num==16'd1567) begin
		isPrime = 1;
	end	else if (num==16'd1571) begin
		isPrime = 1;
	end	else if (num==16'd1579) begin
		isPrime = 1;
	end	else if (num==16'd1583) begin
		isPrime = 1;
	end	else if (num==16'd1597) begin
		isPrime = 1;
	end	else if (num==16'd1601) begin
		isPrime = 1;
	end	else if (num==16'd1607) begin
		isPrime = 1;
	end	else if (num==16'd1609) begin
		isPrime = 1;
	end	else if (num==16'd1613) begin
		isPrime = 1;
	end	else if (num==16'd1619) begin
		isPrime = 1;
	end	else if (num==16'd1621) begin
		isPrime = 1;
	end	else if (num==16'd1627) begin
		isPrime = 1;
	end	else if (num==16'd1637) begin
		isPrime = 1;
	end	else if (num==16'd1657) begin
		isPrime = 1;
	end	else if (num==16'd1663) begin
		isPrime = 1;
	end	else if (num==16'd1667) begin
		isPrime = 1;
	end	else if (num==16'd1669) begin
		isPrime = 1;
	end	else if (num==16'd1693) begin
		isPrime = 1;
	end	else if (num==16'd1697) begin
		isPrime = 1;
	end	else if (num==16'd1699) begin
		isPrime = 1;
	end	else if (num==16'd1709) begin
		isPrime = 1;
	end	else if (num==16'd1721) begin
		isPrime = 1;
	end	else if (num==16'd1723) begin
		isPrime = 1;
	end	else if (num==16'd1733) begin
		isPrime = 1;
	end	else if (num==16'd1741) begin
		isPrime = 1;
	end	else if (num==16'd1747) begin
		isPrime = 1;
	end	else if (num==16'd1753) begin
		isPrime = 1;
	end	else if (num==16'd1759) begin
		isPrime = 1;
	end	else if (num==16'd1777) begin
		isPrime = 1;
	end	else if (num==16'd1783) begin
		isPrime = 1;
	end	else if (num==16'd1787) begin
		isPrime = 1;
	end	else if (num==16'd1789) begin
		isPrime = 1;
	end	else if (num==16'd1801) begin
		isPrime = 1;
	end	else if (num==16'd1811) begin
		isPrime = 1;
	end	else if (num==16'd1823) begin
		isPrime = 1;
	end	else if (num==16'd1831) begin
		isPrime = 1;
	end	else if (num==16'd1847) begin
		isPrime = 1;
	end	else if (num==16'd1861) begin
		isPrime = 1;
	end	else if (num==16'd1867) begin
		isPrime = 1;
	end	else if (num==16'd1871) begin
		isPrime = 1;
	end	else if (num==16'd1873) begin
		isPrime = 1;
	end	else if (num==16'd1877) begin
		isPrime = 1;
	end	else if (num==16'd1879) begin
		isPrime = 1;
	end	else if (num==16'd1889) begin
		isPrime = 1;
	end	else if (num==16'd1901) begin
		isPrime = 1;
	end	else if (num==16'd1907) begin
		isPrime = 1;
	end	else if (num==16'd1913) begin
		isPrime = 1;
	end	else if (num==16'd1931) begin
		isPrime = 1;
	end	else if (num==16'd1933) begin
		isPrime = 1;
	end	else if (num==16'd1949) begin
		isPrime = 1;
	end	else if (num==16'd1951) begin
		isPrime = 1;
	end	else if (num==16'd1973) begin
		isPrime = 1;
	end	else if (num==16'd1979) begin
		isPrime = 1;
	end	else if (num==16'd1987) begin
		isPrime = 1;
	end	else if (num==16'd1993) begin
		isPrime = 1;
	end	else if (num==16'd1997) begin
		isPrime = 1;
	end	else if (num==16'd1999) begin
		isPrime = 1;
	end	else if (num==16'd2003) begin
		isPrime = 1;
	end	else if (num==16'd2011) begin
		isPrime = 1;
	end	else if (num==16'd2017) begin
		isPrime = 1;
	end	else if (num==16'd2027) begin
		isPrime = 1;
	end	else if (num==16'd2029) begin
		isPrime = 1;
	end	else if (num==16'd2039) begin
		isPrime = 1;
	end	else if (num==16'd2053) begin
		isPrime = 1;
	end	else if (num==16'd2063) begin
		isPrime = 1;
	end	else if (num==16'd2069) begin
		isPrime = 1;
	end	else if (num==16'd2081) begin
		isPrime = 1;
	end	else if (num==16'd2083) begin
		isPrime = 1;
	end	else if (num==16'd2087) begin
		isPrime = 1;
	end	else if (num==16'd2089) begin
		isPrime = 1;
	end	else if (num==16'd2099) begin
		isPrime = 1;
	end	else if (num==16'd2111) begin
		isPrime = 1;
	end	else if (num==16'd2113) begin
		isPrime = 1;
	end	else if (num==16'd2129) begin
		isPrime = 1;
	end	else if (num==16'd2131) begin
		isPrime = 1;
	end	else if (num==16'd2137) begin
		isPrime = 1;
	end	else if (num==16'd2141) begin
		isPrime = 1;
	end	else if (num==16'd2143) begin
		isPrime = 1;
	end	else if (num==16'd2153) begin
		isPrime = 1;
	end	else if (num==16'd2161) begin
		isPrime = 1;
	end	else if (num==16'd2179) begin
		isPrime = 1;
	end	else if (num==16'd2203) begin
		isPrime = 1;
	end	else if (num==16'd2207) begin
		isPrime = 1;
	end	else if (num==16'd2213) begin
		isPrime = 1;
	end	else if (num==16'd2221) begin
		isPrime = 1;
	end	else if (num==16'd2237) begin
		isPrime = 1;
	end	else if (num==16'd2239) begin
		isPrime = 1;
	end	else if (num==16'd2243) begin
		isPrime = 1;
	end	else if (num==16'd2251) begin
		isPrime = 1;
	end	else if (num==16'd2267) begin
		isPrime = 1;
	end	else if (num==16'd2269) begin
		isPrime = 1;
	end	else if (num==16'd2273) begin
		isPrime = 1;
	end	else if (num==16'd2281) begin
		isPrime = 1;
	end	else if (num==16'd2287) begin
		isPrime = 1;
	end	else if (num==16'd2293) begin
		isPrime = 1;
	end	else if (num==16'd2297) begin
		isPrime = 1;
	end	else if (num==16'd2309) begin
		isPrime = 1;
	end	else if (num==16'd2311) begin
		isPrime = 1;
	end	else if (num==16'd2333) begin
		isPrime = 1;
	end	else if (num==16'd2339) begin
		isPrime = 1;
	end	else if (num==16'd2341) begin
		isPrime = 1;
	end	else if (num==16'd2347) begin
		isPrime = 1;
	end	else if (num==16'd2351) begin
		isPrime = 1;
	end	else if (num==16'd2357) begin
		isPrime = 1;
	end	else if (num==16'd2371) begin
		isPrime = 1;
	end	else if (num==16'd2377) begin
		isPrime = 1;
	end	else if (num==16'd2381) begin
		isPrime = 1;
	end	else if (num==16'd2383) begin
		isPrime = 1;
	end	else if (num==16'd2389) begin
		isPrime = 1;
	end	else if (num==16'd2393) begin
		isPrime = 1;
	end	else if (num==16'd2399) begin
		isPrime = 1;
	end	else if (num==16'd2411) begin
		isPrime = 1;
	end	else if (num==16'd2417) begin
		isPrime = 1;
	end	else if (num==16'd2423) begin
		isPrime = 1;
	end	else if (num==16'd2437) begin
		isPrime = 1;
	end	else if (num==16'd2441) begin
		isPrime = 1;
	end	else if (num==16'd2447) begin
		isPrime = 1;
	end	else if (num==16'd2459) begin
		isPrime = 1;
	end	else if (num==16'd2467) begin
		isPrime = 1;
	end	else if (num==16'd2473) begin
		isPrime = 1;
	end	else if (num==16'd2477) begin
		isPrime = 1;
	end	else if (num==16'd2503) begin
		isPrime = 1;
	end	else if (num==16'd2521) begin
		isPrime = 1;
	end	else if (num==16'd2531) begin
		isPrime = 1;
	end	else if (num==16'd2539) begin
		isPrime = 1;
	end	else if (num==16'd2543) begin
		isPrime = 1;
	end	else if (num==16'd2549) begin
		isPrime = 1;
	end	else if (num==16'd2551) begin
		isPrime = 1;
	end	else if (num==16'd2557) begin
		isPrime = 1;
	end	else if (num==16'd2579) begin
		isPrime = 1;
	end	else if (num==16'd2591) begin
		isPrime = 1;
	end	else if (num==16'd2593) begin
		isPrime = 1;
	end	else if (num==16'd2609) begin
		isPrime = 1;
	end	else if (num==16'd2617) begin
		isPrime = 1;
	end	else if (num==16'd2621) begin
		isPrime = 1;
	end	else if (num==16'd2633) begin
		isPrime = 1;
	end	else if (num==16'd2647) begin
		isPrime = 1;
	end	else if (num==16'd2657) begin
		isPrime = 1;
	end	else if (num==16'd2659) begin
		isPrime = 1;
	end	else if (num==16'd2663) begin
		isPrime = 1;
	end	else if (num==16'd2671) begin
		isPrime = 1;
	end	else if (num==16'd2677) begin
		isPrime = 1;
	end	else if (num==16'd2683) begin
		isPrime = 1;
	end	else if (num==16'd2687) begin
		isPrime = 1;
	end	else if (num==16'd2689) begin
		isPrime = 1;
	end	else if (num==16'd2693) begin
		isPrime = 1;
	end	else if (num==16'd2699) begin
		isPrime = 1;
	end	else if (num==16'd2707) begin
		isPrime = 1;
	end	else if (num==16'd2711) begin
		isPrime = 1;
	end	else if (num==16'd2713) begin
		isPrime = 1;
	end	else if (num==16'd2719) begin
		isPrime = 1;
	end	else if (num==16'd2729) begin
		isPrime = 1;
	end	else if (num==16'd2731) begin
		isPrime = 1;
	end	else if (num==16'd2741) begin
		isPrime = 1;
	end	else if (num==16'd2749) begin
		isPrime = 1;
	end	else if (num==16'd2753) begin
		isPrime = 1;
	end	else if (num==16'd2767) begin
		isPrime = 1;
	end	else if (num==16'd2777) begin
		isPrime = 1;
	end	else if (num==16'd2789) begin
		isPrime = 1;
	end	else if (num==16'd2791) begin
		isPrime = 1;
	end	else if (num==16'd2797) begin
		isPrime = 1;
	end	else if (num==16'd2801) begin
		isPrime = 1;
	end	else if (num==16'd2803) begin
		isPrime = 1;
	end	else if (num==16'd2819) begin
		isPrime = 1;
	end	else if (num==16'd2833) begin
		isPrime = 1;
	end	else if (num==16'd2837) begin
		isPrime = 1;
	end	else if (num==16'd2843) begin
		isPrime = 1;
	end	else if (num==16'd2851) begin
		isPrime = 1;
	end	else if (num==16'd2857) begin
		isPrime = 1;
	end	else if (num==16'd2861) begin
		isPrime = 1;
	end	else if (num==16'd2879) begin
		isPrime = 1;
	end	else if (num==16'd2887) begin
		isPrime = 1;
	end	else if (num==16'd2897) begin
		isPrime = 1;
	end	else if (num==16'd2903) begin
		isPrime = 1;
	end	else if (num==16'd2909) begin
		isPrime = 1;
	end	else if (num==16'd2917) begin
		isPrime = 1;
	end	else if (num==16'd2927) begin
		isPrime = 1;
	end	else if (num==16'd2939) begin
		isPrime = 1;
	end	else if (num==16'd2953) begin
		isPrime = 1;
	end	else if (num==16'd2957) begin
		isPrime = 1;
	end	else if (num==16'd2963) begin
		isPrime = 1;
	end	else if (num==16'd2969) begin
		isPrime = 1;
	end	else if (num==16'd2971) begin
		isPrime = 1;
	end	else if (num==16'd2999) begin
		isPrime = 1;
	end	else if (num==16'd3001) begin
		isPrime = 1;
	end	else if (num==16'd3011) begin
		isPrime = 1;
	end	else if (num==16'd3019) begin
		isPrime = 1;
	end	else if (num==16'd3023) begin
		isPrime = 1;
	end	else if (num==16'd3037) begin
		isPrime = 1;
	end	else if (num==16'd3041) begin
		isPrime = 1;
	end	else if (num==16'd3049) begin
		isPrime = 1;
	end	else if (num==16'd3061) begin
		isPrime = 1;
	end	else if (num==16'd3067) begin
		isPrime = 1;
	end	else if (num==16'd3079) begin
		isPrime = 1;
	end	else if (num==16'd3083) begin
		isPrime = 1;
	end	else if (num==16'd3089) begin
		isPrime = 1;
	end	else if (num==16'd3109) begin
		isPrime = 1;
	end	else if (num==16'd3119) begin
		isPrime = 1;
	end	else if (num==16'd3121) begin
		isPrime = 1;
	end	else if (num==16'd3137) begin
		isPrime = 1;
	end	else if (num==16'd3163) begin
		isPrime = 1;
	end	else if (num==16'd3167) begin
		isPrime = 1;
	end	else if (num==16'd3169) begin
		isPrime = 1;
	end	else if (num==16'd3181) begin
		isPrime = 1;
	end	else if (num==16'd3187) begin
		isPrime = 1;
	end	else if (num==16'd3191) begin
		isPrime = 1;
	end	else if (num==16'd3203) begin
		isPrime = 1;
	end	else if (num==16'd3209) begin
		isPrime = 1;
	end	else if (num==16'd3217) begin
		isPrime = 1;
	end	else if (num==16'd3221) begin
		isPrime = 1;
	end	else if (num==16'd3229) begin
		isPrime = 1;
	end	else if (num==16'd3251) begin
		isPrime = 1;
	end	else if (num==16'd3253) begin
		isPrime = 1;
	end	else if (num==16'd3257) begin
		isPrime = 1;
	end	else if (num==16'd3259) begin
		isPrime = 1;
	end	else if (num==16'd3271) begin
		isPrime = 1;
	end	else if (num==16'd3299) begin
		isPrime = 1;
	end	else if (num==16'd3301) begin
		isPrime = 1;
	end	else if (num==16'd3307) begin
		isPrime = 1;
	end	else if (num==16'd3313) begin
		isPrime = 1;
	end	else if (num==16'd3319) begin
		isPrime = 1;
	end	else if (num==16'd3323) begin
		isPrime = 1;
	end	else if (num==16'd3329) begin
		isPrime = 1;
	end	else if (num==16'd3331) begin
		isPrime = 1;
	end	else if (num==16'd3343) begin
		isPrime = 1;
	end	else if (num==16'd3347) begin
		isPrime = 1;
	end	else if (num==16'd3359) begin
		isPrime = 1;
	end	else if (num==16'd3361) begin
		isPrime = 1;
	end	else if (num==16'd3371) begin
		isPrime = 1;
	end	else if (num==16'd3373) begin
		isPrime = 1;
	end	else if (num==16'd3389) begin
		isPrime = 1;
	end	else if (num==16'd3391) begin
		isPrime = 1;
	end	else if (num==16'd3407) begin
		isPrime = 1;
	end	else if (num==16'd3413) begin
		isPrime = 1;
	end	else if (num==16'd3433) begin
		isPrime = 1;
	end	else if (num==16'd3449) begin
		isPrime = 1;
	end	else if (num==16'd3457) begin
		isPrime = 1;
	end	else if (num==16'd3461) begin
		isPrime = 1;
	end	else if (num==16'd3463) begin
		isPrime = 1;
	end	else if (num==16'd3467) begin
		isPrime = 1;
	end	else if (num==16'd3469) begin
		isPrime = 1;
	end	else if (num==16'd3491) begin
		isPrime = 1;
	end	else if (num==16'd3499) begin
		isPrime = 1;
	end	else if (num==16'd3511) begin
		isPrime = 1;
	end	else if (num==16'd3517) begin
		isPrime = 1;
	end	else if (num==16'd3527) begin
		isPrime = 1;
	end	else if (num==16'd3529) begin
		isPrime = 1;
	end	else if (num==16'd3533) begin
		isPrime = 1;
	end	else if (num==16'd3539) begin
		isPrime = 1;
	end	else if (num==16'd3541) begin
		isPrime = 1;
	end	else if (num==16'd3547) begin
		isPrime = 1;
	end	else if (num==16'd3557) begin
		isPrime = 1;
	end	else if (num==16'd3559) begin
		isPrime = 1;
	end	else if (num==16'd3571) begin
		isPrime = 1;
	end	else if (num==16'd3581) begin
		isPrime = 1;
	end	else if (num==16'd3583) begin
		isPrime = 1;
	end	else if (num==16'd3593) begin
		isPrime = 1;
	end	else if (num==16'd3607) begin
		isPrime = 1;
	end	else if (num==16'd3613) begin
		isPrime = 1;
	end	else if (num==16'd3617) begin
		isPrime = 1;
	end	else if (num==16'd3623) begin
		isPrime = 1;
	end	else if (num==16'd3631) begin
		isPrime = 1;
	end	else if (num==16'd3637) begin
		isPrime = 1;
	end	else if (num==16'd3643) begin
		isPrime = 1;
	end	else if (num==16'd3659) begin
		isPrime = 1;
	end	else if (num==16'd3671) begin
		isPrime = 1;
	end	else if (num==16'd3673) begin
		isPrime = 1;
	end	else if (num==16'd3677) begin
		isPrime = 1;
	end	else if (num==16'd3691) begin
		isPrime = 1;
	end	else if (num==16'd3697) begin
		isPrime = 1;
	end	else if (num==16'd3701) begin
		isPrime = 1;
	end	else if (num==16'd3709) begin
		isPrime = 1;
	end	else if (num==16'd3719) begin
		isPrime = 1;
	end	else if (num==16'd3727) begin
		isPrime = 1;
	end	else if (num==16'd3733) begin
		isPrime = 1;
	end	else if (num==16'd3739) begin
		isPrime = 1;
	end	else if (num==16'd3761) begin
		isPrime = 1;
	end	else if (num==16'd3767) begin
		isPrime = 1;
	end	else if (num==16'd3769) begin
		isPrime = 1;
	end	else if (num==16'd3779) begin
		isPrime = 1;
	end	else if (num==16'd3793) begin
		isPrime = 1;
	end	else if (num==16'd3797) begin
		isPrime = 1;
	end	else if (num==16'd3803) begin
		isPrime = 1;
	end	else if (num==16'd3821) begin
		isPrime = 1;
	end	else if (num==16'd3823) begin
		isPrime = 1;
	end	else if (num==16'd3833) begin
		isPrime = 1;
	end	else if (num==16'd3847) begin
		isPrime = 1;
	end	else if (num==16'd3851) begin
		isPrime = 1;
	end	else if (num==16'd3853) begin
		isPrime = 1;
	end	else if (num==16'd3863) begin
		isPrime = 1;
	end	else if (num==16'd3877) begin
		isPrime = 1;
	end	else if (num==16'd3881) begin
		isPrime = 1;
	end	else if (num==16'd3889) begin
		isPrime = 1;
	end	else if (num==16'd3907) begin
		isPrime = 1;
	end	else if (num==16'd3911) begin
		isPrime = 1;
	end	else if (num==16'd3917) begin
		isPrime = 1;
	end	else if (num==16'd3919) begin
		isPrime = 1;
	end	else if (num==16'd3923) begin
		isPrime = 1;
	end	else if (num==16'd3929) begin
		isPrime = 1;
	end	else if (num==16'd3931) begin
		isPrime = 1;
	end	else if (num==16'd3943) begin
		isPrime = 1;
	end	else if (num==16'd3947) begin
		isPrime = 1;
	end	else if (num==16'd3967) begin
		isPrime = 1;
	end	else if (num==16'd3989) begin
		isPrime = 1;
	end	else if (num==16'd4001) begin
		isPrime = 1;
	end	else if (num==16'd4003) begin
		isPrime = 1;
	end	else if (num==16'd4007) begin
		isPrime = 1;
	end	else if (num==16'd4013) begin
		isPrime = 1;
	end	else if (num==16'd4019) begin
		isPrime = 1;
	end	else if (num==16'd4021) begin
		isPrime = 1;
	end	else if (num==16'd4027) begin
		isPrime = 1;
	end	else if (num==16'd4049) begin
		isPrime = 1;
	end	else if (num==16'd4051) begin
		isPrime = 1;
	end	else if (num==16'd4057) begin
		isPrime = 1;
	end	else if (num==16'd4073) begin
		isPrime = 1;
	end	else if (num==16'd4079) begin
		isPrime = 1;
	end	else if (num==16'd4091) begin
		isPrime = 1;
	end	else if (num==16'd4093) begin
		isPrime = 1;
	end	else if (num==16'd4099) begin
		isPrime = 1;
	end	else if (num==16'd4111) begin
		isPrime = 1;
	end	else if (num==16'd4127) begin
		isPrime = 1;
	end	else if (num==16'd4129) begin
		isPrime = 1;
	end	else if (num==16'd4133) begin
		isPrime = 1;
	end	else if (num==16'd4139) begin
		isPrime = 1;
	end	else if (num==16'd4153) begin
		isPrime = 1;
	end	else if (num==16'd4157) begin
		isPrime = 1;
	end	else if (num==16'd4159) begin
		isPrime = 1;
	end	else if (num==16'd4177) begin
		isPrime = 1;
	end	else if (num==16'd4201) begin
		isPrime = 1;
	end	else if (num==16'd4211) begin
		isPrime = 1;
	end	else if (num==16'd4217) begin
		isPrime = 1;
	end	else if (num==16'd4219) begin
		isPrime = 1;
	end	else if (num==16'd4229) begin
		isPrime = 1;
	end	else if (num==16'd4231) begin
		isPrime = 1;
	end	else if (num==16'd4241) begin
		isPrime = 1;
	end	else if (num==16'd4243) begin
		isPrime = 1;
	end	else if (num==16'd4253) begin
		isPrime = 1;
	end	else if (num==16'd4259) begin
		isPrime = 1;
	end	else if (num==16'd4261) begin
		isPrime = 1;
	end	else if (num==16'd4271) begin
		isPrime = 1;
	end	else if (num==16'd4273) begin
		isPrime = 1;
	end	else if (num==16'd4283) begin
		isPrime = 1;
	end	else if (num==16'd4289) begin
		isPrime = 1;
	end	else if (num==16'd4297) begin
		isPrime = 1;
	end	else if (num==16'd4327) begin
		isPrime = 1;
	end	else if (num==16'd4337) begin
		isPrime = 1;
	end	else if (num==16'd4339) begin
		isPrime = 1;
	end	else if (num==16'd4349) begin
		isPrime = 1;
	end	else if (num==16'd4357) begin
		isPrime = 1;
	end	else if (num==16'd4363) begin
		isPrime = 1;
	end	else if (num==16'd4373) begin
		isPrime = 1;
	end	else if (num==16'd4391) begin
		isPrime = 1;
	end	else if (num==16'd4397) begin
		isPrime = 1;
	end	else if (num==16'd4409) begin
		isPrime = 1;
	end	else if (num==16'd4421) begin
		isPrime = 1;
	end	else if (num==16'd4423) begin
		isPrime = 1;
	end	else if (num==16'd4441) begin
		isPrime = 1;
	end	else if (num==16'd4447) begin
		isPrime = 1;
	end	else if (num==16'd4451) begin
		isPrime = 1;
	end	else if (num==16'd4457) begin
		isPrime = 1;
	end	else if (num==16'd4463) begin
		isPrime = 1;
	end	else if (num==16'd4481) begin
		isPrime = 1;
	end	else if (num==16'd4483) begin
		isPrime = 1;
	end	else if (num==16'd4493) begin
		isPrime = 1;
	end	else if (num==16'd4507) begin
		isPrime = 1;
	end	else if (num==16'd4513) begin
		isPrime = 1;
	end	else if (num==16'd4517) begin
		isPrime = 1;
	end	else if (num==16'd4519) begin
		isPrime = 1;
	end	else if (num==16'd4523) begin
		isPrime = 1;
	end	else if (num==16'd4547) begin
		isPrime = 1;
	end	else if (num==16'd4549) begin
		isPrime = 1;
	end	else if (num==16'd4561) begin
		isPrime = 1;
	end	else if (num==16'd4567) begin
		isPrime = 1;
	end	else if (num==16'd4583) begin
		isPrime = 1;
	end	else if (num==16'd4591) begin
		isPrime = 1;
	end	else if (num==16'd4597) begin
		isPrime = 1;
	end	else if (num==16'd4603) begin
		isPrime = 1;
	end	else if (num==16'd4621) begin
		isPrime = 1;
	end	else if (num==16'd4637) begin
		isPrime = 1;
	end	else if (num==16'd4639) begin
		isPrime = 1;
	end	else if (num==16'd4643) begin
		isPrime = 1;
	end	else if (num==16'd4649) begin
		isPrime = 1;
	end	else if (num==16'd4651) begin
		isPrime = 1;
	end	else if (num==16'd4657) begin
		isPrime = 1;
	end	else if (num==16'd4663) begin
		isPrime = 1;
	end	else if (num==16'd4673) begin
		isPrime = 1;
	end	else if (num==16'd4679) begin
		isPrime = 1;
	end	else if (num==16'd4691) begin
		isPrime = 1;
	end	else if (num==16'd4703) begin
		isPrime = 1;
	end	else if (num==16'd4721) begin
		isPrime = 1;
	end	else if (num==16'd4723) begin
		isPrime = 1;
	end	else if (num==16'd4729) begin
		isPrime = 1;
	end	else if (num==16'd4733) begin
		isPrime = 1;
	end	else if (num==16'd4751) begin
		isPrime = 1;
	end	else if (num==16'd4759) begin
		isPrime = 1;
	end	else if (num==16'd4783) begin
		isPrime = 1;
	end	else if (num==16'd4787) begin
		isPrime = 1;
	end	else if (num==16'd4789) begin
		isPrime = 1;
	end	else if (num==16'd4793) begin
		isPrime = 1;
	end	else if (num==16'd4799) begin
		isPrime = 1;
	end	else if (num==16'd4801) begin
		isPrime = 1;
	end	else if (num==16'd4813) begin
		isPrime = 1;
	end	else if (num==16'd4817) begin
		isPrime = 1;
	end	else if (num==16'd4831) begin
		isPrime = 1;
	end	else if (num==16'd4861) begin
		isPrime = 1;
	end	else if (num==16'd4871) begin
		isPrime = 1;
	end	else if (num==16'd4877) begin
		isPrime = 1;
	end	else if (num==16'd4889) begin
		isPrime = 1;
	end	else if (num==16'd4903) begin
		isPrime = 1;
	end	else if (num==16'd4909) begin
		isPrime = 1;
	end	else if (num==16'd4919) begin
		isPrime = 1;
	end	else if (num==16'd4931) begin
		isPrime = 1;
	end	else if (num==16'd4933) begin
		isPrime = 1;
	end	else if (num==16'd4937) begin
		isPrime = 1;
	end	else if (num==16'd4943) begin
		isPrime = 1;
	end	else if (num==16'd4951) begin
		isPrime = 1;
	end	else if (num==16'd4957) begin
		isPrime = 1;
	end	else if (num==16'd4967) begin
		isPrime = 1;
	end	else if (num==16'd4969) begin
		isPrime = 1;
	end	else if (num==16'd4973) begin
		isPrime = 1;
	end	else if (num==16'd4987) begin
		isPrime = 1;
	end	else if (num==16'd4993) begin
		isPrime = 1;
	end	else if (num==16'd4999) begin
		isPrime = 1;
	end	else if (num==16'd5003) begin
		isPrime = 1;
	end	else if (num==16'd5009) begin
		isPrime = 1;
	end	else if (num==16'd5011) begin
		isPrime = 1;
	end	else if (num==16'd5021) begin
		isPrime = 1;
	end	else if (num==16'd5023) begin
		isPrime = 1;
	end	else if (num==16'd5039) begin
		isPrime = 1;
	end	else if (num==16'd5051) begin
		isPrime = 1;
	end	else if (num==16'd5059) begin
		isPrime = 1;
	end	else if (num==16'd5077) begin
		isPrime = 1;
	end	else if (num==16'd5081) begin
		isPrime = 1;
	end	else if (num==16'd5087) begin
		isPrime = 1;
	end	else if (num==16'd5099) begin
		isPrime = 1;
	end	else if (num==16'd5101) begin
		isPrime = 1;
	end	else if (num==16'd5107) begin
		isPrime = 1;
	end	else if (num==16'd5113) begin
		isPrime = 1;
	end	else if (num==16'd5119) begin
		isPrime = 1;
	end	else if (num==16'd5147) begin
		isPrime = 1;
	end	else if (num==16'd5153) begin
		isPrime = 1;
	end	else if (num==16'd5167) begin
		isPrime = 1;
	end	else if (num==16'd5171) begin
		isPrime = 1;
	end	else if (num==16'd5179) begin
		isPrime = 1;
	end	else if (num==16'd5189) begin
		isPrime = 1;
	end	else if (num==16'd5197) begin
		isPrime = 1;
	end	else if (num==16'd5209) begin
		isPrime = 1;
	end	else if (num==16'd5227) begin
		isPrime = 1;
	end	else if (num==16'd5231) begin
		isPrime = 1;
	end	else if (num==16'd5233) begin
		isPrime = 1;
	end	else if (num==16'd5237) begin
		isPrime = 1;
	end	else if (num==16'd5261) begin
		isPrime = 1;
	end	else if (num==16'd5273) begin
		isPrime = 1;
	end	else if (num==16'd5279) begin
		isPrime = 1;
	end	else if (num==16'd5281) begin
		isPrime = 1;
	end	else if (num==16'd5297) begin
		isPrime = 1;
	end	else if (num==16'd5303) begin
		isPrime = 1;
	end	else if (num==16'd5309) begin
		isPrime = 1;
	end	else if (num==16'd5323) begin
		isPrime = 1;
	end	else if (num==16'd5333) begin
		isPrime = 1;
	end	else if (num==16'd5347) begin
		isPrime = 1;
	end	else if (num==16'd5351) begin
		isPrime = 1;
	end	else if (num==16'd5381) begin
		isPrime = 1;
	end	else if (num==16'd5387) begin
		isPrime = 1;
	end	else if (num==16'd5393) begin
		isPrime = 1;
	end	else if (num==16'd5399) begin
		isPrime = 1;
	end	else if (num==16'd5407) begin
		isPrime = 1;
	end	else if (num==16'd5413) begin
		isPrime = 1;
	end	else if (num==16'd5417) begin
		isPrime = 1;
	end	else if (num==16'd5419) begin
		isPrime = 1;
	end	else if (num==16'd5431) begin
		isPrime = 1;
	end	else if (num==16'd5437) begin
		isPrime = 1;
	end	else if (num==16'd5441) begin
		isPrime = 1;
	end	else if (num==16'd5443) begin
		isPrime = 1;
	end	else if (num==16'd5449) begin
		isPrime = 1;
	end	else if (num==16'd5471) begin
		isPrime = 1;
	end	else if (num==16'd5477) begin
		isPrime = 1;
	end	else if (num==16'd5479) begin
		isPrime = 1;
	end	else if (num==16'd5483) begin
		isPrime = 1;
	end	else if (num==16'd5501) begin
		isPrime = 1;
	end	else if (num==16'd5503) begin
		isPrime = 1;
	end	else if (num==16'd5507) begin
		isPrime = 1;
	end	else if (num==16'd5519) begin
		isPrime = 1;
	end	else if (num==16'd5521) begin
		isPrime = 1;
	end	else if (num==16'd5527) begin
		isPrime = 1;
	end	else if (num==16'd5531) begin
		isPrime = 1;
	end	else if (num==16'd5557) begin
		isPrime = 1;
	end	else if (num==16'd5563) begin
		isPrime = 1;
	end	else if (num==16'd5569) begin
		isPrime = 1;
	end	else if (num==16'd5573) begin
		isPrime = 1;
	end	else if (num==16'd5581) begin
		isPrime = 1;
	end	else if (num==16'd5591) begin
		isPrime = 1;
	end	else if (num==16'd5623) begin
		isPrime = 1;
	end	else if (num==16'd5639) begin
		isPrime = 1;
	end	else if (num==16'd5641) begin
		isPrime = 1;
	end	else if (num==16'd5647) begin
		isPrime = 1;
	end	else if (num==16'd5651) begin
		isPrime = 1;
	end	else if (num==16'd5653) begin
		isPrime = 1;
	end	else if (num==16'd5657) begin
		isPrime = 1;
	end	else if (num==16'd5659) begin
		isPrime = 1;
	end	else if (num==16'd5669) begin
		isPrime = 1;
	end	else if (num==16'd5683) begin
		isPrime = 1;
	end	else if (num==16'd5689) begin
		isPrime = 1;
	end	else if (num==16'd5693) begin
		isPrime = 1;
	end	else if (num==16'd5701) begin
		isPrime = 1;
	end	else if (num==16'd5711) begin
		isPrime = 1;
	end	else if (num==16'd5717) begin
		isPrime = 1;
	end	else if (num==16'd5737) begin
		isPrime = 1;
	end	else if (num==16'd5741) begin
		isPrime = 1;
	end	else if (num==16'd5743) begin
		isPrime = 1;
	end	else if (num==16'd5749) begin
		isPrime = 1;
	end	else if (num==16'd5779) begin
		isPrime = 1;
	end	else if (num==16'd5783) begin
		isPrime = 1;
	end	else if (num==16'd5791) begin
		isPrime = 1;
	end	else if (num==16'd5801) begin
		isPrime = 1;
	end	else if (num==16'd5807) begin
		isPrime = 1;
	end	else if (num==16'd5813) begin
		isPrime = 1;
	end	else if (num==16'd5821) begin
		isPrime = 1;
	end	else if (num==16'd5827) begin
		isPrime = 1;
	end	else if (num==16'd5839) begin
		isPrime = 1;
	end	else if (num==16'd5843) begin
		isPrime = 1;
	end	else if (num==16'd5849) begin
		isPrime = 1;
	end	else if (num==16'd5851) begin
		isPrime = 1;
	end	else if (num==16'd5857) begin
		isPrime = 1;
	end	else if (num==16'd5861) begin
		isPrime = 1;
	end	else if (num==16'd5867) begin
		isPrime = 1;
	end	else if (num==16'd5869) begin
		isPrime = 1;
	end	else if (num==16'd5879) begin
		isPrime = 1;
	end	else if (num==16'd5881) begin
		isPrime = 1;
	end	else if (num==16'd5897) begin
		isPrime = 1;
	end	else if (num==16'd5903) begin
		isPrime = 1;
	end	else if (num==16'd5923) begin
		isPrime = 1;
	end	else if (num==16'd5927) begin
		isPrime = 1;
	end	else if (num==16'd5939) begin
		isPrime = 1;
	end	else if (num==16'd5953) begin
		isPrime = 1;
	end	else if (num==16'd5981) begin
		isPrime = 1;
	end	else if (num==16'd5987) begin
		isPrime = 1;
	end	else if (num==16'd6007) begin
		isPrime = 1;
	end	else if (num==16'd6011) begin
		isPrime = 1;
	end	else if (num==16'd6029) begin
		isPrime = 1;
	end	else if (num==16'd6037) begin
		isPrime = 1;
	end	else if (num==16'd6043) begin
		isPrime = 1;
	end	else if (num==16'd6047) begin
		isPrime = 1;
	end	else if (num==16'd6053) begin
		isPrime = 1;
	end	else if (num==16'd6067) begin
		isPrime = 1;
	end	else if (num==16'd6073) begin
		isPrime = 1;
	end	else if (num==16'd6079) begin
		isPrime = 1;
	end	else if (num==16'd6089) begin
		isPrime = 1;
	end	else if (num==16'd6091) begin
		isPrime = 1;
	end	else if (num==16'd6101) begin
		isPrime = 1;
	end	else if (num==16'd6113) begin
		isPrime = 1;
	end	else if (num==16'd6121) begin
		isPrime = 1;
	end	else if (num==16'd6131) begin
		isPrime = 1;
	end	else if (num==16'd6133) begin
		isPrime = 1;
	end	else if (num==16'd6143) begin
		isPrime = 1;
	end	else if (num==16'd6151) begin
		isPrime = 1;
	end	else if (num==16'd6163) begin
		isPrime = 1;
	end	else if (num==16'd6173) begin
		isPrime = 1;
	end	else if (num==16'd6197) begin
		isPrime = 1;
	end	else if (num==16'd6199) begin
		isPrime = 1;
	end	else if (num==16'd6203) begin
		isPrime = 1;
	end	else if (num==16'd6211) begin
		isPrime = 1;
	end	else if (num==16'd6217) begin
		isPrime = 1;
	end	else if (num==16'd6221) begin
		isPrime = 1;
	end	else if (num==16'd6229) begin
		isPrime = 1;
	end	else if (num==16'd6247) begin
		isPrime = 1;
	end	else if (num==16'd6257) begin
		isPrime = 1;
	end	else if (num==16'd6263) begin
		isPrime = 1;
	end	else if (num==16'd6269) begin
		isPrime = 1;
	end	else if (num==16'd6271) begin
		isPrime = 1;
	end	else if (num==16'd6277) begin
		isPrime = 1;
	end	else if (num==16'd6287) begin
		isPrime = 1;
	end	else if (num==16'd6299) begin
		isPrime = 1;
	end	else if (num==16'd6301) begin
		isPrime = 1;
	end	else if (num==16'd6311) begin
		isPrime = 1;
	end	else if (num==16'd6317) begin
		isPrime = 1;
	end	else if (num==16'd6323) begin
		isPrime = 1;
	end	else if (num==16'd6329) begin
		isPrime = 1;
	end	else if (num==16'd6337) begin
		isPrime = 1;
	end	else if (num==16'd6343) begin
		isPrime = 1;
	end	else if (num==16'd6353) begin
		isPrime = 1;
	end	else if (num==16'd6359) begin
		isPrime = 1;
	end	else if (num==16'd6361) begin
		isPrime = 1;
	end	else if (num==16'd6367) begin
		isPrime = 1;
	end	else if (num==16'd6373) begin
		isPrime = 1;
	end	else if (num==16'd6379) begin
		isPrime = 1;
	end	else if (num==16'd6389) begin
		isPrime = 1;
	end	else if (num==16'd6397) begin
		isPrime = 1;
	end	else if (num==16'd6421) begin
		isPrime = 1;
	end	else if (num==16'd6427) begin
		isPrime = 1;
	end	else if (num==16'd6449) begin
		isPrime = 1;
	end	else if (num==16'd6451) begin
		isPrime = 1;
	end	else if (num==16'd6469) begin
		isPrime = 1;
	end	else if (num==16'd6473) begin
		isPrime = 1;
	end	else if (num==16'd6481) begin
		isPrime = 1;
	end	else if (num==16'd6491) begin
		isPrime = 1;
	end	else if (num==16'd6521) begin
		isPrime = 1;
	end	else if (num==16'd6529) begin
		isPrime = 1;
	end	else if (num==16'd6547) begin
		isPrime = 1;
	end	else if (num==16'd6551) begin
		isPrime = 1;
	end	else if (num==16'd6553) begin
		isPrime = 1;
	end	else if (num==16'd6563) begin
		isPrime = 1;
	end	else if (num==16'd6569) begin
		isPrime = 1;
	end	else if (num==16'd6571) begin
		isPrime = 1;
	end	else if (num==16'd6577) begin
		isPrime = 1;
	end	else if (num==16'd6581) begin
		isPrime = 1;
	end	else if (num==16'd6599) begin
		isPrime = 1;
	end	else if (num==16'd6607) begin
		isPrime = 1;
	end	else if (num==16'd6619) begin
		isPrime = 1;
	end	else if (num==16'd6637) begin
		isPrime = 1;
	end	else if (num==16'd6653) begin
		isPrime = 1;
	end	else if (num==16'd6659) begin
		isPrime = 1;
	end	else if (num==16'd6661) begin
		isPrime = 1;
	end	else if (num==16'd6673) begin
		isPrime = 1;
	end	else if (num==16'd6679) begin
		isPrime = 1;
	end	else if (num==16'd6689) begin
		isPrime = 1;
	end	else if (num==16'd6691) begin
		isPrime = 1;
	end	else if (num==16'd6701) begin
		isPrime = 1;
	end	else if (num==16'd6703) begin
		isPrime = 1;
	end	else if (num==16'd6709) begin
		isPrime = 1;
	end	else if (num==16'd6719) begin
		isPrime = 1;
	end	else if (num==16'd6733) begin
		isPrime = 1;
	end	else if (num==16'd6737) begin
		isPrime = 1;
	end	else if (num==16'd6761) begin
		isPrime = 1;
	end	else if (num==16'd6763) begin
		isPrime = 1;
	end	else if (num==16'd6779) begin
		isPrime = 1;
	end	else if (num==16'd6781) begin
		isPrime = 1;
	end	else if (num==16'd6791) begin
		isPrime = 1;
	end	else if (num==16'd6793) begin
		isPrime = 1;
	end	else if (num==16'd6803) begin
		isPrime = 1;
	end	else if (num==16'd6823) begin
		isPrime = 1;
	end	else if (num==16'd6827) begin
		isPrime = 1;
	end	else if (num==16'd6829) begin
		isPrime = 1;
	end	else if (num==16'd6833) begin
		isPrime = 1;
	end	else if (num==16'd6841) begin
		isPrime = 1;
	end	else if (num==16'd6857) begin
		isPrime = 1;
	end	else if (num==16'd6863) begin
		isPrime = 1;
	end	else if (num==16'd6869) begin
		isPrime = 1;
	end	else if (num==16'd6871) begin
		isPrime = 1;
	end	else if (num==16'd6883) begin
		isPrime = 1;
	end	else if (num==16'd6899) begin
		isPrime = 1;
	end	else if (num==16'd6907) begin
		isPrime = 1;
	end	else if (num==16'd6911) begin
		isPrime = 1;
	end	else if (num==16'd6917) begin
		isPrime = 1;
	end	else if (num==16'd6947) begin
		isPrime = 1;
	end	else if (num==16'd6949) begin
		isPrime = 1;
	end	else if (num==16'd6959) begin
		isPrime = 1;
	end	else if (num==16'd6961) begin
		isPrime = 1;
	end	else if (num==16'd6967) begin
		isPrime = 1;
	end	else if (num==16'd6971) begin
		isPrime = 1;
	end	else if (num==16'd6977) begin
		isPrime = 1;
	end	else if (num==16'd6983) begin
		isPrime = 1;
	end	else if (num==16'd6991) begin
		isPrime = 1;
	end	else if (num==16'd6997) begin
		isPrime = 1;
	end	else if (num==16'd7001) begin
		isPrime = 1;
	end	else if (num==16'd7013) begin
		isPrime = 1;
	end	else if (num==16'd7019) begin
		isPrime = 1;
	end	else if (num==16'd7027) begin
		isPrime = 1;
	end	else if (num==16'd7039) begin
		isPrime = 1;
	end	else if (num==16'd7043) begin
		isPrime = 1;
	end	else if (num==16'd7057) begin
		isPrime = 1;
	end	else if (num==16'd7069) begin
		isPrime = 1;
	end	else if (num==16'd7079) begin
		isPrime = 1;
	end	else if (num==16'd7103) begin
		isPrime = 1;
	end	else if (num==16'd7109) begin
		isPrime = 1;
	end	else if (num==16'd7121) begin
		isPrime = 1;
	end	else if (num==16'd7127) begin
		isPrime = 1;
	end	else if (num==16'd7129) begin
		isPrime = 1;
	end	else if (num==16'd7151) begin
		isPrime = 1;
	end	else if (num==16'd7159) begin
		isPrime = 1;
	end	else if (num==16'd7177) begin
		isPrime = 1;
	end	else if (num==16'd7187) begin
		isPrime = 1;
	end	else if (num==16'd7193) begin
		isPrime = 1;
	end	else if (num==16'd7207) begin
		isPrime = 1;
	end	else if (num==16'd7211) begin
		isPrime = 1;
	end	else if (num==16'd7213) begin
		isPrime = 1;
	end	else if (num==16'd7219) begin
		isPrime = 1;
	end	else if (num==16'd7229) begin
		isPrime = 1;
	end	else if (num==16'd7237) begin
		isPrime = 1;
	end	else if (num==16'd7243) begin
		isPrime = 1;
	end	else if (num==16'd7247) begin
		isPrime = 1;
	end	else if (num==16'd7253) begin
		isPrime = 1;
	end	else if (num==16'd7283) begin
		isPrime = 1;
	end	else if (num==16'd7297) begin
		isPrime = 1;
	end	else if (num==16'd7307) begin
		isPrime = 1;
	end	else if (num==16'd7309) begin
		isPrime = 1;
	end	else if (num==16'd7321) begin
		isPrime = 1;
	end	else if (num==16'd7331) begin
		isPrime = 1;
	end	else if (num==16'd7333) begin
		isPrime = 1;
	end	else if (num==16'd7349) begin
		isPrime = 1;
	end	else if (num==16'd7351) begin
		isPrime = 1;
	end	else if (num==16'd7369) begin
		isPrime = 1;
	end	else if (num==16'd7393) begin
		isPrime = 1;
	end	else if (num==16'd7411) begin
		isPrime = 1;
	end	else if (num==16'd7417) begin
		isPrime = 1;
	end	else if (num==16'd7433) begin
		isPrime = 1;
	end	else if (num==16'd7451) begin
		isPrime = 1;
	end	else if (num==16'd7457) begin
		isPrime = 1;
	end	else if (num==16'd7459) begin
		isPrime = 1;
	end	else if (num==16'd7477) begin
		isPrime = 1;
	end	else if (num==16'd7481) begin
		isPrime = 1;
	end	else if (num==16'd7487) begin
		isPrime = 1;
	end	else if (num==16'd7489) begin
		isPrime = 1;
	end	else if (num==16'd7499) begin
		isPrime = 1;
	end	else if (num==16'd7507) begin
		isPrime = 1;
	end	else if (num==16'd7517) begin
		isPrime = 1;
	end	else if (num==16'd7523) begin
		isPrime = 1;
	end	else if (num==16'd7529) begin
		isPrime = 1;
	end	else if (num==16'd7537) begin
		isPrime = 1;
	end	else if (num==16'd7541) begin
		isPrime = 1;
	end	else if (num==16'd7547) begin
		isPrime = 1;
	end	else if (num==16'd7549) begin
		isPrime = 1;
	end	else if (num==16'd7559) begin
		isPrime = 1;
	end	else if (num==16'd7561) begin
		isPrime = 1;
	end	else if (num==16'd7573) begin
		isPrime = 1;
	end	else if (num==16'd7577) begin
		isPrime = 1;
	end	else if (num==16'd7583) begin
		isPrime = 1;
	end	else if (num==16'd7589) begin
		isPrime = 1;
	end	else if (num==16'd7591) begin
		isPrime = 1;
	end	else if (num==16'd7603) begin
		isPrime = 1;
	end	else if (num==16'd7607) begin
		isPrime = 1;
	end	else if (num==16'd7621) begin
		isPrime = 1;
	end	else if (num==16'd7639) begin
		isPrime = 1;
	end	else if (num==16'd7643) begin
		isPrime = 1;
	end	else if (num==16'd7649) begin
		isPrime = 1;
	end	else if (num==16'd7669) begin
		isPrime = 1;
	end	else if (num==16'd7673) begin
		isPrime = 1;
	end	else if (num==16'd7681) begin
		isPrime = 1;
	end	else if (num==16'd7687) begin
		isPrime = 1;
	end	else if (num==16'd7691) begin
		isPrime = 1;
	end	else if (num==16'd7699) begin
		isPrime = 1;
	end	else if (num==16'd7703) begin
		isPrime = 1;
	end	else if (num==16'd7717) begin
		isPrime = 1;
	end	else if (num==16'd7723) begin
		isPrime = 1;
	end	else if (num==16'd7727) begin
		isPrime = 1;
	end	else if (num==16'd7741) begin
		isPrime = 1;
	end	else if (num==16'd7753) begin
		isPrime = 1;
	end	else if (num==16'd7757) begin
		isPrime = 1;
	end	else if (num==16'd7759) begin
		isPrime = 1;
	end	else if (num==16'd7789) begin
		isPrime = 1;
	end	else if (num==16'd7793) begin
		isPrime = 1;
	end	else if (num==16'd7817) begin
		isPrime = 1;
	end	else if (num==16'd7823) begin
		isPrime = 1;
	end	else if (num==16'd7829) begin
		isPrime = 1;
	end	else if (num==16'd7841) begin
		isPrime = 1;
	end	else if (num==16'd7853) begin
		isPrime = 1;
	end	else if (num==16'd7867) begin
		isPrime = 1;
	end	else if (num==16'd7873) begin
		isPrime = 1;
	end	else if (num==16'd7877) begin
		isPrime = 1;
	end	else if (num==16'd7879) begin
		isPrime = 1;
	end	else if (num==16'd7883) begin
		isPrime = 1;
	end	else if (num==16'd7901) begin
		isPrime = 1;
	end	else if (num==16'd7907) begin
		isPrime = 1;
	end	else if (num==16'd7919) begin
		isPrime = 1;
	end	else if (num==16'd7927) begin
		isPrime = 1;
	end	else if (num==16'd7933) begin
		isPrime = 1;
	end	else if (num==16'd7937) begin
		isPrime = 1;
	end	else if (num==16'd7949) begin
		isPrime = 1;
	end	else if (num==16'd7951) begin
		isPrime = 1;
	end	else if (num==16'd7963) begin
		isPrime = 1;
	end	else if (num==16'd7993) begin
		isPrime = 1;
	end	else if (num==16'd8009) begin
		isPrime = 1;
	end	else if (num==16'd8011) begin
		isPrime = 1;
	end	else if (num==16'd8017) begin
		isPrime = 1;
	end	else if (num==16'd8039) begin
		isPrime = 1;
	end	else if (num==16'd8053) begin
		isPrime = 1;
	end	else if (num==16'd8059) begin
		isPrime = 1;
	end	else if (num==16'd8069) begin
		isPrime = 1;
	end	else if (num==16'd8081) begin
		isPrime = 1;
	end	else if (num==16'd8087) begin
		isPrime = 1;
	end	else if (num==16'd8089) begin
		isPrime = 1;
	end	else if (num==16'd8093) begin
		isPrime = 1;
	end	else if (num==16'd8101) begin
		isPrime = 1;
	end	else if (num==16'd8111) begin
		isPrime = 1;
	end	else if (num==16'd8117) begin
		isPrime = 1;
	end	else if (num==16'd8123) begin
		isPrime = 1;
	end	else if (num==16'd8147) begin
		isPrime = 1;
	end	else if (num==16'd8161) begin
		isPrime = 1;
	end	else if (num==16'd8167) begin
		isPrime = 1;
	end	else if (num==16'd8171) begin
		isPrime = 1;
	end	else if (num==16'd8179) begin
		isPrime = 1;
	end	else if (num==16'd8191) begin
		isPrime = 1;
	end	else if (num==16'd8209) begin
		isPrime = 1;
	end	else if (num==16'd8219) begin
		isPrime = 1;
	end	else if (num==16'd8221) begin
		isPrime = 1;
	end	else if (num==16'd8231) begin
		isPrime = 1;
	end	else if (num==16'd8233) begin
		isPrime = 1;
	end	else if (num==16'd8237) begin
		isPrime = 1;
	end	else if (num==16'd8243) begin
		isPrime = 1;
	end	else if (num==16'd8263) begin
		isPrime = 1;
	end	else if (num==16'd8269) begin
		isPrime = 1;
	end	else if (num==16'd8273) begin
		isPrime = 1;
	end	else if (num==16'd8287) begin
		isPrime = 1;
	end	else if (num==16'd8291) begin
		isPrime = 1;
	end	else if (num==16'd8293) begin
		isPrime = 1;
	end	else if (num==16'd8297) begin
		isPrime = 1;
	end	else if (num==16'd8311) begin
		isPrime = 1;
	end	else if (num==16'd8317) begin
		isPrime = 1;
	end	else if (num==16'd8329) begin
		isPrime = 1;
	end	else if (num==16'd8353) begin
		isPrime = 1;
	end	else if (num==16'd8363) begin
		isPrime = 1;
	end	else if (num==16'd8369) begin
		isPrime = 1;
	end	else if (num==16'd8377) begin
		isPrime = 1;
	end	else if (num==16'd8387) begin
		isPrime = 1;
	end	else if (num==16'd8389) begin
		isPrime = 1;
	end	else if (num==16'd8419) begin
		isPrime = 1;
	end	else if (num==16'd8423) begin
		isPrime = 1;
	end	else if (num==16'd8429) begin
		isPrime = 1;
	end	else if (num==16'd8431) begin
		isPrime = 1;
	end	else if (num==16'd8443) begin
		isPrime = 1;
	end	else if (num==16'd8447) begin
		isPrime = 1;
	end	else if (num==16'd8461) begin
		isPrime = 1;
	end	else if (num==16'd8467) begin
		isPrime = 1;
	end	else if (num==16'd8501) begin
		isPrime = 1;
	end	else if (num==16'd8513) begin
		isPrime = 1;
	end	else if (num==16'd8521) begin
		isPrime = 1;
	end	else if (num==16'd8527) begin
		isPrime = 1;
	end	else if (num==16'd8537) begin
		isPrime = 1;
	end	else if (num==16'd8539) begin
		isPrime = 1;
	end	else if (num==16'd8543) begin
		isPrime = 1;
	end	else if (num==16'd8563) begin
		isPrime = 1;
	end	else if (num==16'd8573) begin
		isPrime = 1;
	end	else if (num==16'd8581) begin
		isPrime = 1;
	end	else if (num==16'd8597) begin
		isPrime = 1;
	end	else if (num==16'd8599) begin
		isPrime = 1;
	end	else if (num==16'd8609) begin
		isPrime = 1;
	end	else if (num==16'd8623) begin
		isPrime = 1;
	end	else if (num==16'd8627) begin
		isPrime = 1;
	end	else if (num==16'd8629) begin
		isPrime = 1;
	end	else if (num==16'd8641) begin
		isPrime = 1;
	end	else if (num==16'd8647) begin
		isPrime = 1;
	end	else if (num==16'd8663) begin
		isPrime = 1;
	end	else if (num==16'd8669) begin
		isPrime = 1;
	end	else if (num==16'd8677) begin
		isPrime = 1;
	end	else if (num==16'd8681) begin
		isPrime = 1;
	end	else if (num==16'd8689) begin
		isPrime = 1;
	end	else if (num==16'd8693) begin
		isPrime = 1;
	end	else if (num==16'd8699) begin
		isPrime = 1;
	end	else if (num==16'd8707) begin
		isPrime = 1;
	end	else if (num==16'd8713) begin
		isPrime = 1;
	end	else if (num==16'd8719) begin
		isPrime = 1;
	end	else if (num==16'd8731) begin
		isPrime = 1;
	end	else if (num==16'd8737) begin
		isPrime = 1;
	end	else if (num==16'd8741) begin
		isPrime = 1;
	end	else if (num==16'd8747) begin
		isPrime = 1;
	end	else if (num==16'd8753) begin
		isPrime = 1;
	end	else if (num==16'd8761) begin
		isPrime = 1;
	end	else if (num==16'd8779) begin
		isPrime = 1;
	end	else if (num==16'd8783) begin
		isPrime = 1;
	end	else if (num==16'd8803) begin
		isPrime = 1;
	end	else if (num==16'd8807) begin
		isPrime = 1;
	end	else if (num==16'd8819) begin
		isPrime = 1;
	end	else if (num==16'd8821) begin
		isPrime = 1;
	end	else if (num==16'd8831) begin
		isPrime = 1;
	end	else if (num==16'd8837) begin
		isPrime = 1;
	end	else if (num==16'd8839) begin
		isPrime = 1;
	end	else if (num==16'd8849) begin
		isPrime = 1;
	end	else if (num==16'd8861) begin
		isPrime = 1;
	end	else if (num==16'd8863) begin
		isPrime = 1;
	end	else if (num==16'd8867) begin
		isPrime = 1;
	end	else if (num==16'd8887) begin
		isPrime = 1;
	end	else if (num==16'd8893) begin
		isPrime = 1;
	end	else if (num==16'd8923) begin
		isPrime = 1;
	end	else if (num==16'd8929) begin
		isPrime = 1;
	end	else if (num==16'd8933) begin
		isPrime = 1;
	end	else if (num==16'd8941) begin
		isPrime = 1;
	end	else if (num==16'd8951) begin
		isPrime = 1;
	end	else if (num==16'd8963) begin
		isPrime = 1;
	end	else if (num==16'd8969) begin
		isPrime = 1;
	end	else if (num==16'd8971) begin
		isPrime = 1;
	end	else if (num==16'd8999) begin
		isPrime = 1;
	end	else if (num==16'd9001) begin
		isPrime = 1;
	end	else if (num==16'd9007) begin
		isPrime = 1;
	end	else if (num==16'd9011) begin
		isPrime = 1;
	end	else if (num==16'd9013) begin
		isPrime = 1;
	end	else if (num==16'd9029) begin
		isPrime = 1;
	end	else if (num==16'd9041) begin
		isPrime = 1;
	end	else if (num==16'd9043) begin
		isPrime = 1;
	end	else if (num==16'd9049) begin
		isPrime = 1;
	end	else if (num==16'd9059) begin
		isPrime = 1;
	end	else if (num==16'd9067) begin
		isPrime = 1;
	end	else if (num==16'd9091) begin
		isPrime = 1;
	end	else if (num==16'd9103) begin
		isPrime = 1;
	end	else if (num==16'd9109) begin
		isPrime = 1;
	end	else if (num==16'd9127) begin
		isPrime = 1;
	end	else if (num==16'd9133) begin
		isPrime = 1;
	end	else if (num==16'd9137) begin
		isPrime = 1;
	end	else if (num==16'd9151) begin
		isPrime = 1;
	end	else if (num==16'd9157) begin
		isPrime = 1;
	end	else if (num==16'd9161) begin
		isPrime = 1;
	end	else if (num==16'd9173) begin
		isPrime = 1;
	end	else if (num==16'd9181) begin
		isPrime = 1;
	end	else if (num==16'd9187) begin
		isPrime = 1;
	end	else if (num==16'd9199) begin
		isPrime = 1;
	end	else if (num==16'd9203) begin
		isPrime = 1;
	end	else if (num==16'd9209) begin
		isPrime = 1;
	end	else if (num==16'd9221) begin
		isPrime = 1;
	end	else if (num==16'd9227) begin
		isPrime = 1;
	end	else if (num==16'd9239) begin
		isPrime = 1;
	end	else if (num==16'd9241) begin
		isPrime = 1;
	end	else if (num==16'd9257) begin
		isPrime = 1;
	end	else if (num==16'd9277) begin
		isPrime = 1;
	end	else if (num==16'd9281) begin
		isPrime = 1;
	end	else if (num==16'd9283) begin
		isPrime = 1;
	end	else if (num==16'd9293) begin
		isPrime = 1;
	end	else if (num==16'd9311) begin
		isPrime = 1;
	end	else if (num==16'd9319) begin
		isPrime = 1;
	end	else if (num==16'd9323) begin
		isPrime = 1;
	end	else if (num==16'd9337) begin
		isPrime = 1;
	end	else if (num==16'd9341) begin
		isPrime = 1;
	end	else if (num==16'd9343) begin
		isPrime = 1;
	end	else if (num==16'd9349) begin
		isPrime = 1;
	end	else if (num==16'd9371) begin
		isPrime = 1;
	end	else if (num==16'd9377) begin
		isPrime = 1;
	end	else if (num==16'd9391) begin
		isPrime = 1;
	end	else if (num==16'd9397) begin
		isPrime = 1;
	end	else if (num==16'd9403) begin
		isPrime = 1;
	end	else if (num==16'd9413) begin
		isPrime = 1;
	end	else if (num==16'd9419) begin
		isPrime = 1;
	end	else if (num==16'd9421) begin
		isPrime = 1;
	end	else if (num==16'd9431) begin
		isPrime = 1;
	end	else if (num==16'd9433) begin
		isPrime = 1;
	end	else if (num==16'd9437) begin
		isPrime = 1;
	end	else if (num==16'd9439) begin
		isPrime = 1;
	end	else if (num==16'd9461) begin
		isPrime = 1;
	end	else if (num==16'd9463) begin
		isPrime = 1;
	end	else if (num==16'd9467) begin
		isPrime = 1;
	end	else if (num==16'd9473) begin
		isPrime = 1;
	end	else if (num==16'd9479) begin
		isPrime = 1;
	end	else if (num==16'd9491) begin
		isPrime = 1;
	end	else if (num==16'd9497) begin
		isPrime = 1;
	end	else if (num==16'd9511) begin
		isPrime = 1;
	end	else if (num==16'd9521) begin
		isPrime = 1;
	end	else if (num==16'd9533) begin
		isPrime = 1;
	end	else if (num==16'd9539) begin
		isPrime = 1;
	end	else if (num==16'd9547) begin
		isPrime = 1;
	end	else if (num==16'd9551) begin
		isPrime = 1;
	end	else if (num==16'd9587) begin
		isPrime = 1;
	end	else if (num==16'd9601) begin
		isPrime = 1;
	end	else if (num==16'd9613) begin
		isPrime = 1;
	end	else if (num==16'd9619) begin
		isPrime = 1;
	end	else if (num==16'd9623) begin
		isPrime = 1;
	end	else if (num==16'd9629) begin
		isPrime = 1;
	end	else if (num==16'd9631) begin
		isPrime = 1;
	end	else if (num==16'd9643) begin
		isPrime = 1;
	end	else if (num==16'd9649) begin
		isPrime = 1;
	end	else if (num==16'd9661) begin
		isPrime = 1;
	end	else if (num==16'd9677) begin
		isPrime = 1;
	end	else if (num==16'd9679) begin
		isPrime = 1;
	end	else if (num==16'd9689) begin
		isPrime = 1;
	end	else if (num==16'd9697) begin
		isPrime = 1;
	end	else if (num==16'd9719) begin
		isPrime = 1;
	end	else if (num==16'd9721) begin
		isPrime = 1;
	end	else if (num==16'd9733) begin
		isPrime = 1;
	end	else if (num==16'd9739) begin
		isPrime = 1;
	end	else if (num==16'd9743) begin
		isPrime = 1;
	end	else if (num==16'd9749) begin
		isPrime = 1;
	end	else if (num==16'd9767) begin
		isPrime = 1;
	end	else if (num==16'd9769) begin
		isPrime = 1;
	end	else if (num==16'd9781) begin
		isPrime = 1;
	end	else if (num==16'd9787) begin
		isPrime = 1;
	end	else if (num==16'd9791) begin
		isPrime = 1;
	end	else if (num==16'd9803) begin
		isPrime = 1;
	end	else if (num==16'd9811) begin
		isPrime = 1;
	end	else if (num==16'd9817) begin
		isPrime = 1;
	end	else if (num==16'd9829) begin
		isPrime = 1;
	end	else if (num==16'd9833) begin
		isPrime = 1;
	end	else if (num==16'd9839) begin
		isPrime = 1;
	end	else if (num==16'd9851) begin
		isPrime = 1;
	end	else if (num==16'd9857) begin
		isPrime = 1;
	end	else if (num==16'd9859) begin
		isPrime = 1;
	end	else if (num==16'd9871) begin
		isPrime = 1;
	end	else if (num==16'd9883) begin
		isPrime = 1;
	end	else if (num==16'd9887) begin
		isPrime = 1;
	end	else if (num==16'd9901) begin
		isPrime = 1;
	end	else if (num==16'd9907) begin
		isPrime = 1;
	end	else if (num==16'd9923) begin
		isPrime = 1;
	end	else if (num==16'd9929) begin
		isPrime = 1;
	end	else if (num==16'd9931) begin
		isPrime = 1;
	end	else if (num==16'd9941) begin
		isPrime = 1;
	end	else if (num==16'd9949) begin
		isPrime = 1;
	end	else if (num==16'd9967) begin
		isPrime = 1;
	end	else if (num==16'd9973) begin
		isPrime = 1;
	end	else if (num==16'd10007) begin
		isPrime = 1;
	end	else if (num==16'd10009) begin
		isPrime = 1;
	end	else if (num==16'd10037) begin
		isPrime = 1;
	end	else if (num==16'd10039) begin
		isPrime = 1;
	end	else if (num==16'd10061) begin
		isPrime = 1;
	end	else if (num==16'd10067) begin
		isPrime = 1;
	end	else if (num==16'd10069) begin
		isPrime = 1;
	end	else if (num==16'd10079) begin
		isPrime = 1;
	end	else if (num==16'd10091) begin
		isPrime = 1;
	end	else if (num==16'd10093) begin
		isPrime = 1;
	end	else if (num==16'd10099) begin
		isPrime = 1;
	end	else if (num==16'd10103) begin
		isPrime = 1;
	end	else if (num==16'd10111) begin
		isPrime = 1;
	end	else if (num==16'd10133) begin
		isPrime = 1;
	end	else if (num==16'd10139) begin
		isPrime = 1;
	end	else if (num==16'd10141) begin
		isPrime = 1;
	end	else if (num==16'd10151) begin
		isPrime = 1;
	end	else if (num==16'd10159) begin
		isPrime = 1;
	end	else if (num==16'd10163) begin
		isPrime = 1;
	end	else if (num==16'd10169) begin
		isPrime = 1;
	end	else if (num==16'd10177) begin
		isPrime = 1;
	end	else if (num==16'd10181) begin
		isPrime = 1;
	end	else if (num==16'd10193) begin
		isPrime = 1;
	end	else if (num==16'd10211) begin
		isPrime = 1;
	end	else if (num==16'd10223) begin
		isPrime = 1;
	end	else if (num==16'd10243) begin
		isPrime = 1;
	end	else if (num==16'd10247) begin
		isPrime = 1;
	end	else if (num==16'd10253) begin
		isPrime = 1;
	end	else if (num==16'd10259) begin
		isPrime = 1;
	end	else if (num==16'd10267) begin
		isPrime = 1;
	end	else if (num==16'd10271) begin
		isPrime = 1;
	end	else if (num==16'd10273) begin
		isPrime = 1;
	end	else if (num==16'd10289) begin
		isPrime = 1;
	end	else if (num==16'd10301) begin
		isPrime = 1;
	end	else if (num==16'd10303) begin
		isPrime = 1;
	end	else if (num==16'd10313) begin
		isPrime = 1;
	end	else if (num==16'd10321) begin
		isPrime = 1;
	end	else if (num==16'd10331) begin
		isPrime = 1;
	end	else if (num==16'd10333) begin
		isPrime = 1;
	end	else if (num==16'd10337) begin
		isPrime = 1;
	end	else if (num==16'd10343) begin
		isPrime = 1;
	end	else if (num==16'd10357) begin
		isPrime = 1;
	end	else if (num==16'd10369) begin
		isPrime = 1;
	end	else if (num==16'd10391) begin
		isPrime = 1;
	end	else if (num==16'd10399) begin
		isPrime = 1;
	end	else if (num==16'd10427) begin
		isPrime = 1;
	end	else if (num==16'd10429) begin
		isPrime = 1;
	end	else if (num==16'd10433) begin
		isPrime = 1;
	end	else if (num==16'd10453) begin
		isPrime = 1;
	end	else if (num==16'd10457) begin
		isPrime = 1;
	end	else if (num==16'd10459) begin
		isPrime = 1;
	end	else if (num==16'd10463) begin
		isPrime = 1;
	end	else if (num==16'd10477) begin
		isPrime = 1;
	end	else if (num==16'd10487) begin
		isPrime = 1;
	end	else if (num==16'd10499) begin
		isPrime = 1;
	end	else if (num==16'd10501) begin
		isPrime = 1;
	end	else if (num==16'd10513) begin
		isPrime = 1;
	end	else if (num==16'd10529) begin
		isPrime = 1;
	end	else if (num==16'd10531) begin
		isPrime = 1;
	end	else if (num==16'd10559) begin
		isPrime = 1;
	end	else if (num==16'd10567) begin
		isPrime = 1;
	end	else if (num==16'd10589) begin
		isPrime = 1;
	end	else if (num==16'd10597) begin
		isPrime = 1;
	end	else if (num==16'd10601) begin
		isPrime = 1;
	end	else if (num==16'd10607) begin
		isPrime = 1;
	end	else if (num==16'd10613) begin
		isPrime = 1;
	end	else if (num==16'd10627) begin
		isPrime = 1;
	end	else if (num==16'd10631) begin
		isPrime = 1;
	end	else if (num==16'd10639) begin
		isPrime = 1;
	end	else if (num==16'd10651) begin
		isPrime = 1;
	end	else if (num==16'd10657) begin
		isPrime = 1;
	end	else if (num==16'd10663) begin
		isPrime = 1;
	end	else if (num==16'd10667) begin
		isPrime = 1;
	end	else if (num==16'd10687) begin
		isPrime = 1;
	end	else if (num==16'd10691) begin
		isPrime = 1;
	end	else if (num==16'd10709) begin
		isPrime = 1;
	end	else if (num==16'd10711) begin
		isPrime = 1;
	end	else if (num==16'd10723) begin
		isPrime = 1;
	end	else if (num==16'd10729) begin
		isPrime = 1;
	end	else if (num==16'd10733) begin
		isPrime = 1;
	end	else if (num==16'd10739) begin
		isPrime = 1;
	end	else if (num==16'd10753) begin
		isPrime = 1;
	end	else if (num==16'd10771) begin
		isPrime = 1;
	end	else if (num==16'd10781) begin
		isPrime = 1;
	end	else if (num==16'd10789) begin
		isPrime = 1;
	end	else if (num==16'd10799) begin
		isPrime = 1;
	end	else if (num==16'd10831) begin
		isPrime = 1;
	end	else if (num==16'd10837) begin
		isPrime = 1;
	end	else if (num==16'd10847) begin
		isPrime = 1;
	end	else if (num==16'd10853) begin
		isPrime = 1;
	end	else if (num==16'd10859) begin
		isPrime = 1;
	end	else if (num==16'd10861) begin
		isPrime = 1;
	end	else if (num==16'd10867) begin
		isPrime = 1;
	end	else if (num==16'd10883) begin
		isPrime = 1;
	end	else if (num==16'd10889) begin
		isPrime = 1;
	end	else if (num==16'd10891) begin
		isPrime = 1;
	end	else if (num==16'd10903) begin
		isPrime = 1;
	end	else if (num==16'd10909) begin
		isPrime = 1;
	end	else if (num==16'd10937) begin
		isPrime = 1;
	end	else if (num==16'd10939) begin
		isPrime = 1;
	end	else if (num==16'd10949) begin
		isPrime = 1;
	end	else if (num==16'd10957) begin
		isPrime = 1;
	end	else if (num==16'd10973) begin
		isPrime = 1;
	end	else if (num==16'd10979) begin
		isPrime = 1;
	end	else if (num==16'd10987) begin
		isPrime = 1;
	end	else if (num==16'd10993) begin
		isPrime = 1;
	end	else if (num==16'd11003) begin
		isPrime = 1;
	end	else if (num==16'd11027) begin
		isPrime = 1;
	end	else if (num==16'd11047) begin
		isPrime = 1;
	end	else if (num==16'd11057) begin
		isPrime = 1;
	end	else if (num==16'd11059) begin
		isPrime = 1;
	end	else if (num==16'd11069) begin
		isPrime = 1;
	end	else if (num==16'd11071) begin
		isPrime = 1;
	end	else if (num==16'd11083) begin
		isPrime = 1;
	end	else if (num==16'd11087) begin
		isPrime = 1;
	end	else if (num==16'd11093) begin
		isPrime = 1;
	end	else if (num==16'd11113) begin
		isPrime = 1;
	end	else if (num==16'd11117) begin
		isPrime = 1;
	end	else if (num==16'd11119) begin
		isPrime = 1;
	end	else if (num==16'd11131) begin
		isPrime = 1;
	end	else if (num==16'd11149) begin
		isPrime = 1;
	end	else if (num==16'd11159) begin
		isPrime = 1;
	end	else if (num==16'd11161) begin
		isPrime = 1;
	end	else if (num==16'd11171) begin
		isPrime = 1;
	end	else if (num==16'd11173) begin
		isPrime = 1;
	end	else if (num==16'd11177) begin
		isPrime = 1;
	end	else if (num==16'd11197) begin
		isPrime = 1;
	end	else if (num==16'd11213) begin
		isPrime = 1;
	end	else if (num==16'd11239) begin
		isPrime = 1;
	end	else if (num==16'd11243) begin
		isPrime = 1;
	end	else if (num==16'd11251) begin
		isPrime = 1;
	end	else if (num==16'd11257) begin
		isPrime = 1;
	end	else if (num==16'd11261) begin
		isPrime = 1;
	end	else if (num==16'd11273) begin
		isPrime = 1;
	end	else if (num==16'd11279) begin
		isPrime = 1;
	end	else if (num==16'd11287) begin
		isPrime = 1;
	end	else if (num==16'd11299) begin
		isPrime = 1;
	end	else if (num==16'd11311) begin
		isPrime = 1;
	end	else if (num==16'd11317) begin
		isPrime = 1;
	end	else if (num==16'd11321) begin
		isPrime = 1;
	end	else if (num==16'd11329) begin
		isPrime = 1;
	end	else if (num==16'd11351) begin
		isPrime = 1;
	end	else if (num==16'd11353) begin
		isPrime = 1;
	end	else if (num==16'd11369) begin
		isPrime = 1;
	end	else if (num==16'd11383) begin
		isPrime = 1;
	end	else if (num==16'd11393) begin
		isPrime = 1;
	end	else if (num==16'd11399) begin
		isPrime = 1;
	end	else if (num==16'd11411) begin
		isPrime = 1;
	end	else if (num==16'd11423) begin
		isPrime = 1;
	end	else if (num==16'd11437) begin
		isPrime = 1;
	end	else if (num==16'd11443) begin
		isPrime = 1;
	end	else if (num==16'd11447) begin
		isPrime = 1;
	end	else if (num==16'd11467) begin
		isPrime = 1;
	end	else if (num==16'd11471) begin
		isPrime = 1;
	end	else if (num==16'd11483) begin
		isPrime = 1;
	end	else if (num==16'd11489) begin
		isPrime = 1;
	end	else if (num==16'd11491) begin
		isPrime = 1;
	end	else if (num==16'd11497) begin
		isPrime = 1;
	end	else if (num==16'd11503) begin
		isPrime = 1;
	end	else if (num==16'd11519) begin
		isPrime = 1;
	end	else if (num==16'd11527) begin
		isPrime = 1;
	end	else if (num==16'd11549) begin
		isPrime = 1;
	end	else if (num==16'd11551) begin
		isPrime = 1;
	end	else if (num==16'd11579) begin
		isPrime = 1;
	end	else if (num==16'd11587) begin
		isPrime = 1;
	end	else if (num==16'd11593) begin
		isPrime = 1;
	end	else if (num==16'd11597) begin
		isPrime = 1;
	end	else if (num==16'd11617) begin
		isPrime = 1;
	end	else if (num==16'd11621) begin
		isPrime = 1;
	end	else if (num==16'd11633) begin
		isPrime = 1;
	end	else if (num==16'd11657) begin
		isPrime = 1;
	end	else if (num==16'd11677) begin
		isPrime = 1;
	end	else if (num==16'd11681) begin
		isPrime = 1;
	end	else if (num==16'd11689) begin
		isPrime = 1;
	end	else if (num==16'd11699) begin
		isPrime = 1;
	end	else if (num==16'd11701) begin
		isPrime = 1;
	end	else if (num==16'd11717) begin
		isPrime = 1;
	end	else if (num==16'd11719) begin
		isPrime = 1;
	end	else if (num==16'd11731) begin
		isPrime = 1;
	end	else if (num==16'd11743) begin
		isPrime = 1;
	end	else if (num==16'd11777) begin
		isPrime = 1;
	end	else if (num==16'd11779) begin
		isPrime = 1;
	end	else if (num==16'd11783) begin
		isPrime = 1;
	end	else if (num==16'd11789) begin
		isPrime = 1;
	end	else if (num==16'd11801) begin
		isPrime = 1;
	end	else if (num==16'd11807) begin
		isPrime = 1;
	end	else if (num==16'd11813) begin
		isPrime = 1;
	end	else if (num==16'd11821) begin
		isPrime = 1;
	end	else if (num==16'd11827) begin
		isPrime = 1;
	end	else if (num==16'd11831) begin
		isPrime = 1;
	end	else if (num==16'd11833) begin
		isPrime = 1;
	end	else if (num==16'd11839) begin
		isPrime = 1;
	end	else if (num==16'd11863) begin
		isPrime = 1;
	end	else if (num==16'd11867) begin
		isPrime = 1;
	end	else if (num==16'd11887) begin
		isPrime = 1;
	end	else if (num==16'd11897) begin
		isPrime = 1;
	end	else if (num==16'd11903) begin
		isPrime = 1;
	end	else if (num==16'd11909) begin
		isPrime = 1;
	end	else if (num==16'd11923) begin
		isPrime = 1;
	end	else if (num==16'd11927) begin
		isPrime = 1;
	end	else if (num==16'd11933) begin
		isPrime = 1;
	end	else if (num==16'd11939) begin
		isPrime = 1;
	end	else if (num==16'd11941) begin
		isPrime = 1;
	end	else if (num==16'd11953) begin
		isPrime = 1;
	end	else if (num==16'd11959) begin
		isPrime = 1;
	end	else if (num==16'd11969) begin
		isPrime = 1;
	end	else if (num==16'd11971) begin
		isPrime = 1;
	end	else if (num==16'd11981) begin
		isPrime = 1;
	end	else if (num==16'd11987) begin
		isPrime = 1;
	end	else if (num==16'd12007) begin
		isPrime = 1;
	end	else if (num==16'd12011) begin
		isPrime = 1;
	end	else if (num==16'd12037) begin
		isPrime = 1;
	end	else if (num==16'd12041) begin
		isPrime = 1;
	end	else if (num==16'd12043) begin
		isPrime = 1;
	end	else if (num==16'd12049) begin
		isPrime = 1;
	end	else if (num==16'd12071) begin
		isPrime = 1;
	end	else if (num==16'd12073) begin
		isPrime = 1;
	end	else if (num==16'd12097) begin
		isPrime = 1;
	end	else if (num==16'd12101) begin
		isPrime = 1;
	end	else if (num==16'd12107) begin
		isPrime = 1;
	end	else if (num==16'd12109) begin
		isPrime = 1;
	end	else if (num==16'd12113) begin
		isPrime = 1;
	end	else if (num==16'd12119) begin
		isPrime = 1;
	end	else if (num==16'd12143) begin
		isPrime = 1;
	end	else if (num==16'd12149) begin
		isPrime = 1;
	end	else if (num==16'd12157) begin
		isPrime = 1;
	end	else if (num==16'd12161) begin
		isPrime = 1;
	end	else if (num==16'd12163) begin
		isPrime = 1;
	end	else if (num==16'd12197) begin
		isPrime = 1;
	end	else if (num==16'd12203) begin
		isPrime = 1;
	end	else if (num==16'd12211) begin
		isPrime = 1;
	end	else if (num==16'd12227) begin
		isPrime = 1;
	end	else if (num==16'd12239) begin
		isPrime = 1;
	end	else if (num==16'd12241) begin
		isPrime = 1;
	end	else if (num==16'd12251) begin
		isPrime = 1;
	end	else if (num==16'd12253) begin
		isPrime = 1;
	end	else if (num==16'd12263) begin
		isPrime = 1;
	end	else if (num==16'd12269) begin
		isPrime = 1;
	end	else if (num==16'd12277) begin
		isPrime = 1;
	end	else if (num==16'd12281) begin
		isPrime = 1;
	end	else if (num==16'd12289) begin
		isPrime = 1;
	end	else if (num==16'd12301) begin
		isPrime = 1;
	end	else if (num==16'd12323) begin
		isPrime = 1;
	end	else if (num==16'd12329) begin
		isPrime = 1;
	end	else if (num==16'd12343) begin
		isPrime = 1;
	end	else if (num==16'd12347) begin
		isPrime = 1;
	end	else if (num==16'd12373) begin
		isPrime = 1;
	end	else if (num==16'd12377) begin
		isPrime = 1;
	end	else if (num==16'd12379) begin
		isPrime = 1;
	end	else if (num==16'd12391) begin
		isPrime = 1;
	end	else if (num==16'd12401) begin
		isPrime = 1;
	end	else if (num==16'd12409) begin
		isPrime = 1;
	end	else if (num==16'd12413) begin
		isPrime = 1;
	end	else if (num==16'd12421) begin
		isPrime = 1;
	end	else if (num==16'd12433) begin
		isPrime = 1;
	end	else if (num==16'd12437) begin
		isPrime = 1;
	end	else if (num==16'd12451) begin
		isPrime = 1;
	end	else if (num==16'd12457) begin
		isPrime = 1;
	end	else if (num==16'd12473) begin
		isPrime = 1;
	end	else if (num==16'd12479) begin
		isPrime = 1;
	end	else if (num==16'd12487) begin
		isPrime = 1;
	end	else if (num==16'd12491) begin
		isPrime = 1;
	end	else if (num==16'd12497) begin
		isPrime = 1;
	end	else if (num==16'd12503) begin
		isPrime = 1;
	end	else if (num==16'd12511) begin
		isPrime = 1;
	end	else if (num==16'd12517) begin
		isPrime = 1;
	end	else if (num==16'd12527) begin
		isPrime = 1;
	end	else if (num==16'd12539) begin
		isPrime = 1;
	end	else if (num==16'd12541) begin
		isPrime = 1;
	end	else if (num==16'd12547) begin
		isPrime = 1;
	end	else if (num==16'd12553) begin
		isPrime = 1;
	end	else if (num==16'd12569) begin
		isPrime = 1;
	end	else if (num==16'd12577) begin
		isPrime = 1;
	end	else if (num==16'd12583) begin
		isPrime = 1;
	end	else if (num==16'd12589) begin
		isPrime = 1;
	end	else if (num==16'd12601) begin
		isPrime = 1;
	end	else if (num==16'd12611) begin
		isPrime = 1;
	end	else if (num==16'd12613) begin
		isPrime = 1;
	end	else if (num==16'd12619) begin
		isPrime = 1;
	end	else if (num==16'd12637) begin
		isPrime = 1;
	end	else if (num==16'd12641) begin
		isPrime = 1;
	end	else if (num==16'd12647) begin
		isPrime = 1;
	end	else if (num==16'd12653) begin
		isPrime = 1;
	end	else if (num==16'd12659) begin
		isPrime = 1;
	end	else if (num==16'd12671) begin
		isPrime = 1;
	end	else if (num==16'd12689) begin
		isPrime = 1;
	end	else if (num==16'd12697) begin
		isPrime = 1;
	end	else if (num==16'd12703) begin
		isPrime = 1;
	end	else if (num==16'd12713) begin
		isPrime = 1;
	end	else if (num==16'd12721) begin
		isPrime = 1;
	end	else if (num==16'd12739) begin
		isPrime = 1;
	end	else if (num==16'd12743) begin
		isPrime = 1;
	end	else if (num==16'd12757) begin
		isPrime = 1;
	end	else if (num==16'd12763) begin
		isPrime = 1;
	end	else if (num==16'd12781) begin
		isPrime = 1;
	end	else if (num==16'd12791) begin
		isPrime = 1;
	end	else if (num==16'd12799) begin
		isPrime = 1;
	end	else if (num==16'd12809) begin
		isPrime = 1;
	end	else if (num==16'd12821) begin
		isPrime = 1;
	end	else if (num==16'd12823) begin
		isPrime = 1;
	end	else if (num==16'd12829) begin
		isPrime = 1;
	end	else if (num==16'd12841) begin
		isPrime = 1;
	end	else if (num==16'd12853) begin
		isPrime = 1;
	end	else if (num==16'd12889) begin
		isPrime = 1;
	end	else if (num==16'd12893) begin
		isPrime = 1;
	end	else if (num==16'd12899) begin
		isPrime = 1;
	end	else if (num==16'd12907) begin
		isPrime = 1;
	end	else if (num==16'd12911) begin
		isPrime = 1;
	end	else if (num==16'd12917) begin
		isPrime = 1;
	end	else if (num==16'd12919) begin
		isPrime = 1;
	end	else if (num==16'd12923) begin
		isPrime = 1;
	end	else if (num==16'd12941) begin
		isPrime = 1;
	end	else if (num==16'd12953) begin
		isPrime = 1;
	end	else if (num==16'd12959) begin
		isPrime = 1;
	end	else if (num==16'd12967) begin
		isPrime = 1;
	end	else if (num==16'd12973) begin
		isPrime = 1;
	end	else if (num==16'd12979) begin
		isPrime = 1;
	end	else if (num==16'd12983) begin
		isPrime = 1;
	end	else if (num==16'd13001) begin
		isPrime = 1;
	end	else if (num==16'd13003) begin
		isPrime = 1;
	end	else if (num==16'd13007) begin
		isPrime = 1;
	end	else if (num==16'd13009) begin
		isPrime = 1;
	end	else if (num==16'd13033) begin
		isPrime = 1;
	end	else if (num==16'd13037) begin
		isPrime = 1;
	end	else if (num==16'd13043) begin
		isPrime = 1;
	end	else if (num==16'd13049) begin
		isPrime = 1;
	end	else if (num==16'd13063) begin
		isPrime = 1;
	end	else if (num==16'd13093) begin
		isPrime = 1;
	end	else if (num==16'd13099) begin
		isPrime = 1;
	end	else if (num==16'd13103) begin
		isPrime = 1;
	end	else if (num==16'd13109) begin
		isPrime = 1;
	end	else if (num==16'd13121) begin
		isPrime = 1;
	end	else if (num==16'd13127) begin
		isPrime = 1;
	end	else if (num==16'd13147) begin
		isPrime = 1;
	end	else if (num==16'd13151) begin
		isPrime = 1;
	end	else if (num==16'd13159) begin
		isPrime = 1;
	end	else if (num==16'd13163) begin
		isPrime = 1;
	end	else if (num==16'd13171) begin
		isPrime = 1;
	end	else if (num==16'd13177) begin
		isPrime = 1;
	end	else if (num==16'd13183) begin
		isPrime = 1;
	end	else if (num==16'd13187) begin
		isPrime = 1;
	end	else if (num==16'd13217) begin
		isPrime = 1;
	end	else if (num==16'd13219) begin
		isPrime = 1;
	end	else if (num==16'd13229) begin
		isPrime = 1;
	end	else if (num==16'd13241) begin
		isPrime = 1;
	end	else if (num==16'd13249) begin
		isPrime = 1;
	end	else if (num==16'd13259) begin
		isPrime = 1;
	end	else if (num==16'd13267) begin
		isPrime = 1;
	end	else if (num==16'd13291) begin
		isPrime = 1;
	end	else if (num==16'd13297) begin
		isPrime = 1;
	end	else if (num==16'd13309) begin
		isPrime = 1;
	end	else if (num==16'd13313) begin
		isPrime = 1;
	end	else if (num==16'd13327) begin
		isPrime = 1;
	end	else if (num==16'd13331) begin
		isPrime = 1;
	end	else if (num==16'd13337) begin
		isPrime = 1;
	end	else if (num==16'd13339) begin
		isPrime = 1;
	end	else if (num==16'd13367) begin
		isPrime = 1;
	end	else if (num==16'd13381) begin
		isPrime = 1;
	end	else if (num==16'd13397) begin
		isPrime = 1;
	end	else if (num==16'd13399) begin
		isPrime = 1;
	end	else if (num==16'd13411) begin
		isPrime = 1;
	end	else if (num==16'd13417) begin
		isPrime = 1;
	end	else if (num==16'd13421) begin
		isPrime = 1;
	end	else if (num==16'd13441) begin
		isPrime = 1;
	end	else if (num==16'd13451) begin
		isPrime = 1;
	end	else if (num==16'd13457) begin
		isPrime = 1;
	end	else if (num==16'd13463) begin
		isPrime = 1;
	end	else if (num==16'd13469) begin
		isPrime = 1;
	end	else if (num==16'd13477) begin
		isPrime = 1;
	end	else if (num==16'd13487) begin
		isPrime = 1;
	end	else if (num==16'd13499) begin
		isPrime = 1;
	end	else if (num==16'd13513) begin
		isPrime = 1;
	end	else if (num==16'd13523) begin
		isPrime = 1;
	end	else if (num==16'd13537) begin
		isPrime = 1;
	end	else if (num==16'd13553) begin
		isPrime = 1;
	end	else if (num==16'd13567) begin
		isPrime = 1;
	end	else if (num==16'd13577) begin
		isPrime = 1;
	end	else if (num==16'd13591) begin
		isPrime = 1;
	end	else if (num==16'd13597) begin
		isPrime = 1;
	end	else if (num==16'd13613) begin
		isPrime = 1;
	end	else if (num==16'd13619) begin
		isPrime = 1;
	end	else if (num==16'd13627) begin
		isPrime = 1;
	end	else if (num==16'd13633) begin
		isPrime = 1;
	end	else if (num==16'd13649) begin
		isPrime = 1;
	end	else if (num==16'd13669) begin
		isPrime = 1;
	end	else if (num==16'd13679) begin
		isPrime = 1;
	end	else if (num==16'd13681) begin
		isPrime = 1;
	end	else if (num==16'd13687) begin
		isPrime = 1;
	end	else if (num==16'd13691) begin
		isPrime = 1;
	end	else if (num==16'd13693) begin
		isPrime = 1;
	end	else if (num==16'd13697) begin
		isPrime = 1;
	end	else if (num==16'd13709) begin
		isPrime = 1;
	end	else if (num==16'd13711) begin
		isPrime = 1;
	end	else if (num==16'd13721) begin
		isPrime = 1;
	end	else if (num==16'd13723) begin
		isPrime = 1;
	end	else if (num==16'd13729) begin
		isPrime = 1;
	end	else if (num==16'd13751) begin
		isPrime = 1;
	end	else if (num==16'd13757) begin
		isPrime = 1;
	end	else if (num==16'd13759) begin
		isPrime = 1;
	end	else if (num==16'd13763) begin
		isPrime = 1;
	end	else if (num==16'd13781) begin
		isPrime = 1;
	end	else if (num==16'd13789) begin
		isPrime = 1;
	end	else if (num==16'd13799) begin
		isPrime = 1;
	end	else if (num==16'd13807) begin
		isPrime = 1;
	end	else if (num==16'd13829) begin
		isPrime = 1;
	end	else if (num==16'd13831) begin
		isPrime = 1;
	end	else if (num==16'd13841) begin
		isPrime = 1;
	end	else if (num==16'd13859) begin
		isPrime = 1;
	end	else if (num==16'd13873) begin
		isPrime = 1;
	end	else if (num==16'd13877) begin
		isPrime = 1;
	end	else if (num==16'd13879) begin
		isPrime = 1;
	end	else if (num==16'd13883) begin
		isPrime = 1;
	end	else if (num==16'd13901) begin
		isPrime = 1;
	end	else if (num==16'd13903) begin
		isPrime = 1;
	end	else if (num==16'd13907) begin
		isPrime = 1;
	end	else if (num==16'd13913) begin
		isPrime = 1;
	end	else if (num==16'd13921) begin
		isPrime = 1;
	end	else if (num==16'd13931) begin
		isPrime = 1;
	end	else if (num==16'd13933) begin
		isPrime = 1;
	end	else if (num==16'd13963) begin
		isPrime = 1;
	end	else if (num==16'd13967) begin
		isPrime = 1;
	end	else if (num==16'd13997) begin
		isPrime = 1;
	end	else if (num==16'd13999) begin
		isPrime = 1;
	end	else if (num==16'd14009) begin
		isPrime = 1;
	end	else if (num==16'd14011) begin
		isPrime = 1;
	end	else if (num==16'd14029) begin
		isPrime = 1;
	end	else if (num==16'd14033) begin
		isPrime = 1;
	end	else if (num==16'd14051) begin
		isPrime = 1;
	end	else if (num==16'd14057) begin
		isPrime = 1;
	end	else if (num==16'd14071) begin
		isPrime = 1;
	end	else if (num==16'd14081) begin
		isPrime = 1;
	end	else if (num==16'd14083) begin
		isPrime = 1;
	end	else if (num==16'd14087) begin
		isPrime = 1;
	end	else if (num==16'd14107) begin
		isPrime = 1;
	end	else if (num==16'd14143) begin
		isPrime = 1;
	end	else if (num==16'd14149) begin
		isPrime = 1;
	end	else if (num==16'd14153) begin
		isPrime = 1;
	end	else if (num==16'd14159) begin
		isPrime = 1;
	end	else if (num==16'd14173) begin
		isPrime = 1;
	end	else if (num==16'd14177) begin
		isPrime = 1;
	end	else if (num==16'd14197) begin
		isPrime = 1;
	end	else if (num==16'd14207) begin
		isPrime = 1;
	end	else if (num==16'd14221) begin
		isPrime = 1;
	end	else if (num==16'd14243) begin
		isPrime = 1;
	end	else if (num==16'd14249) begin
		isPrime = 1;
	end	else if (num==16'd14251) begin
		isPrime = 1;
	end	else if (num==16'd14281) begin
		isPrime = 1;
	end	else if (num==16'd14293) begin
		isPrime = 1;
	end	else if (num==16'd14303) begin
		isPrime = 1;
	end	else if (num==16'd14321) begin
		isPrime = 1;
	end	else if (num==16'd14323) begin
		isPrime = 1;
	end	else if (num==16'd14327) begin
		isPrime = 1;
	end	else if (num==16'd14341) begin
		isPrime = 1;
	end	else if (num==16'd14347) begin
		isPrime = 1;
	end	else if (num==16'd14369) begin
		isPrime = 1;
	end	else if (num==16'd14387) begin
		isPrime = 1;
	end	else if (num==16'd14389) begin
		isPrime = 1;
	end	else if (num==16'd14401) begin
		isPrime = 1;
	end	else if (num==16'd14407) begin
		isPrime = 1;
	end	else if (num==16'd14411) begin
		isPrime = 1;
	end	else if (num==16'd14419) begin
		isPrime = 1;
	end	else if (num==16'd14423) begin
		isPrime = 1;
	end	else if (num==16'd14431) begin
		isPrime = 1;
	end	else if (num==16'd14437) begin
		isPrime = 1;
	end	else if (num==16'd14447) begin
		isPrime = 1;
	end	else if (num==16'd14449) begin
		isPrime = 1;
	end	else if (num==16'd14461) begin
		isPrime = 1;
	end	else if (num==16'd14479) begin
		isPrime = 1;
	end	else if (num==16'd14489) begin
		isPrime = 1;
	end	else if (num==16'd14503) begin
		isPrime = 1;
	end	else if (num==16'd14519) begin
		isPrime = 1;
	end	else if (num==16'd14533) begin
		isPrime = 1;
	end	else if (num==16'd14537) begin
		isPrime = 1;
	end	else if (num==16'd14543) begin
		isPrime = 1;
	end	else if (num==16'd14549) begin
		isPrime = 1;
	end	else if (num==16'd14551) begin
		isPrime = 1;
	end	else if (num==16'd14557) begin
		isPrime = 1;
	end	else if (num==16'd14561) begin
		isPrime = 1;
	end	else if (num==16'd14563) begin
		isPrime = 1;
	end	else if (num==16'd14591) begin
		isPrime = 1;
	end	else if (num==16'd14593) begin
		isPrime = 1;
	end	else if (num==16'd14621) begin
		isPrime = 1;
	end	else if (num==16'd14627) begin
		isPrime = 1;
	end	else if (num==16'd14629) begin
		isPrime = 1;
	end	else if (num==16'd14633) begin
		isPrime = 1;
	end	else if (num==16'd14639) begin
		isPrime = 1;
	end	else if (num==16'd14653) begin
		isPrime = 1;
	end	else if (num==16'd14657) begin
		isPrime = 1;
	end	else if (num==16'd14669) begin
		isPrime = 1;
	end	else if (num==16'd14683) begin
		isPrime = 1;
	end	else if (num==16'd14699) begin
		isPrime = 1;
	end	else if (num==16'd14713) begin
		isPrime = 1;
	end	else if (num==16'd14717) begin
		isPrime = 1;
	end	else if (num==16'd14723) begin
		isPrime = 1;
	end	else if (num==16'd14731) begin
		isPrime = 1;
	end	else if (num==16'd14737) begin
		isPrime = 1;
	end	else if (num==16'd14741) begin
		isPrime = 1;
	end	else if (num==16'd14747) begin
		isPrime = 1;
	end	else if (num==16'd14753) begin
		isPrime = 1;
	end	else if (num==16'd14759) begin
		isPrime = 1;
	end	else if (num==16'd14767) begin
		isPrime = 1;
	end	else if (num==16'd14771) begin
		isPrime = 1;
	end	else if (num==16'd14779) begin
		isPrime = 1;
	end	else if (num==16'd14783) begin
		isPrime = 1;
	end	else if (num==16'd14797) begin
		isPrime = 1;
	end	else if (num==16'd14813) begin
		isPrime = 1;
	end	else if (num==16'd14821) begin
		isPrime = 1;
	end	else if (num==16'd14827) begin
		isPrime = 1;
	end	else if (num==16'd14831) begin
		isPrime = 1;
	end	else if (num==16'd14843) begin
		isPrime = 1;
	end	else if (num==16'd14851) begin
		isPrime = 1;
	end	else if (num==16'd14867) begin
		isPrime = 1;
	end	else if (num==16'd14869) begin
		isPrime = 1;
	end	else if (num==16'd14879) begin
		isPrime = 1;
	end	else if (num==16'd14887) begin
		isPrime = 1;
	end	else if (num==16'd14891) begin
		isPrime = 1;
	end	else if (num==16'd14897) begin
		isPrime = 1;
	end	else if (num==16'd14923) begin
		isPrime = 1;
	end	else if (num==16'd14929) begin
		isPrime = 1;
	end	else if (num==16'd14939) begin
		isPrime = 1;
	end	else if (num==16'd14947) begin
		isPrime = 1;
	end	else if (num==16'd14951) begin
		isPrime = 1;
	end	else if (num==16'd14957) begin
		isPrime = 1;
	end	else if (num==16'd14969) begin
		isPrime = 1;
	end	else if (num==16'd14983) begin
		isPrime = 1;
	end	else if (num==16'd15013) begin
		isPrime = 1;
	end	else if (num==16'd15017) begin
		isPrime = 1;
	end	else if (num==16'd15031) begin
		isPrime = 1;
	end	else if (num==16'd15053) begin
		isPrime = 1;
	end	else if (num==16'd15061) begin
		isPrime = 1;
	end	else if (num==16'd15073) begin
		isPrime = 1;
	end	else if (num==16'd15077) begin
		isPrime = 1;
	end	else if (num==16'd15083) begin
		isPrime = 1;
	end	else if (num==16'd15091) begin
		isPrime = 1;
	end	else if (num==16'd15101) begin
		isPrime = 1;
	end	else if (num==16'd15107) begin
		isPrime = 1;
	end	else if (num==16'd15121) begin
		isPrime = 1;
	end	else if (num==16'd15131) begin
		isPrime = 1;
	end	else if (num==16'd15137) begin
		isPrime = 1;
	end	else if (num==16'd15139) begin
		isPrime = 1;
	end	else if (num==16'd15149) begin
		isPrime = 1;
	end	else if (num==16'd15161) begin
		isPrime = 1;
	end	else if (num==16'd15173) begin
		isPrime = 1;
	end	else if (num==16'd15187) begin
		isPrime = 1;
	end	else if (num==16'd15193) begin
		isPrime = 1;
	end	else if (num==16'd15199) begin
		isPrime = 1;
	end	else if (num==16'd15217) begin
		isPrime = 1;
	end	else if (num==16'd15227) begin
		isPrime = 1;
	end	else if (num==16'd15233) begin
		isPrime = 1;
	end	else if (num==16'd15241) begin
		isPrime = 1;
	end	else if (num==16'd15259) begin
		isPrime = 1;
	end	else if (num==16'd15263) begin
		isPrime = 1;
	end	else if (num==16'd15269) begin
		isPrime = 1;
	end	else if (num==16'd15271) begin
		isPrime = 1;
	end	else if (num==16'd15277) begin
		isPrime = 1;
	end	else if (num==16'd15287) begin
		isPrime = 1;
	end	else if (num==16'd15289) begin
		isPrime = 1;
	end	else if (num==16'd15299) begin
		isPrime = 1;
	end	else if (num==16'd15307) begin
		isPrime = 1;
	end	else if (num==16'd15313) begin
		isPrime = 1;
	end	else if (num==16'd15319) begin
		isPrime = 1;
	end	else if (num==16'd15329) begin
		isPrime = 1;
	end	else if (num==16'd15331) begin
		isPrime = 1;
	end	else if (num==16'd15349) begin
		isPrime = 1;
	end	else if (num==16'd15359) begin
		isPrime = 1;
	end	else if (num==16'd15361) begin
		isPrime = 1;
	end	else if (num==16'd15373) begin
		isPrime = 1;
	end	else if (num==16'd15377) begin
		isPrime = 1;
	end	else if (num==16'd15383) begin
		isPrime = 1;
	end	else if (num==16'd15391) begin
		isPrime = 1;
	end	else if (num==16'd15401) begin
		isPrime = 1;
	end	else if (num==16'd15413) begin
		isPrime = 1;
	end	else if (num==16'd15427) begin
		isPrime = 1;
	end	else if (num==16'd15439) begin
		isPrime = 1;
	end	else if (num==16'd15443) begin
		isPrime = 1;
	end	else if (num==16'd15451) begin
		isPrime = 1;
	end	else if (num==16'd15461) begin
		isPrime = 1;
	end	else if (num==16'd15467) begin
		isPrime = 1;
	end	else if (num==16'd15473) begin
		isPrime = 1;
	end	else if (num==16'd15493) begin
		isPrime = 1;
	end	else if (num==16'd15497) begin
		isPrime = 1;
	end	else if (num==16'd15511) begin
		isPrime = 1;
	end	else if (num==16'd15527) begin
		isPrime = 1;
	end	else if (num==16'd15541) begin
		isPrime = 1;
	end	else if (num==16'd15551) begin
		isPrime = 1;
	end	else if (num==16'd15559) begin
		isPrime = 1;
	end	else if (num==16'd15569) begin
		isPrime = 1;
	end	else if (num==16'd15581) begin
		isPrime = 1;
	end	else if (num==16'd15583) begin
		isPrime = 1;
	end	else if (num==16'd15601) begin
		isPrime = 1;
	end	else if (num==16'd15607) begin
		isPrime = 1;
	end	else if (num==16'd15619) begin
		isPrime = 1;
	end	else if (num==16'd15629) begin
		isPrime = 1;
	end	else if (num==16'd15641) begin
		isPrime = 1;
	end	else if (num==16'd15643) begin
		isPrime = 1;
	end	else if (num==16'd15647) begin
		isPrime = 1;
	end	else if (num==16'd15649) begin
		isPrime = 1;
	end	else if (num==16'd15661) begin
		isPrime = 1;
	end	else if (num==16'd15667) begin
		isPrime = 1;
	end	else if (num==16'd15671) begin
		isPrime = 1;
	end	else if (num==16'd15679) begin
		isPrime = 1;
	end	else if (num==16'd15683) begin
		isPrime = 1;
	end	else if (num==16'd15727) begin
		isPrime = 1;
	end	else if (num==16'd15731) begin
		isPrime = 1;
	end	else if (num==16'd15733) begin
		isPrime = 1;
	end	else if (num==16'd15737) begin
		isPrime = 1;
	end	else if (num==16'd15739) begin
		isPrime = 1;
	end	else if (num==16'd15749) begin
		isPrime = 1;
	end	else if (num==16'd15761) begin
		isPrime = 1;
	end	else if (num==16'd15767) begin
		isPrime = 1;
	end	else if (num==16'd15773) begin
		isPrime = 1;
	end	else if (num==16'd15787) begin
		isPrime = 1;
	end	else if (num==16'd15791) begin
		isPrime = 1;
	end	else if (num==16'd15797) begin
		isPrime = 1;
	end	else if (num==16'd15803) begin
		isPrime = 1;
	end	else if (num==16'd15809) begin
		isPrime = 1;
	end	else if (num==16'd15817) begin
		isPrime = 1;
	end	else if (num==16'd15823) begin
		isPrime = 1;
	end	else if (num==16'd15859) begin
		isPrime = 1;
	end	else if (num==16'd15877) begin
		isPrime = 1;
	end	else if (num==16'd15881) begin
		isPrime = 1;
	end	else if (num==16'd15887) begin
		isPrime = 1;
	end	else if (num==16'd15889) begin
		isPrime = 1;
	end	else if (num==16'd15901) begin
		isPrime = 1;
	end	else if (num==16'd15907) begin
		isPrime = 1;
	end	else if (num==16'd15913) begin
		isPrime = 1;
	end	else if (num==16'd15919) begin
		isPrime = 1;
	end	else if (num==16'd15923) begin
		isPrime = 1;
	end	else if (num==16'd15937) begin
		isPrime = 1;
	end	else if (num==16'd15959) begin
		isPrime = 1;
	end	else if (num==16'd15971) begin
		isPrime = 1;
	end	else if (num==16'd15973) begin
		isPrime = 1;
	end	else if (num==16'd15991) begin
		isPrime = 1;
	end	else if (num==16'd16001) begin
		isPrime = 1;
	end	else if (num==16'd16007) begin
		isPrime = 1;
	end	else if (num==16'd16033) begin
		isPrime = 1;
	end	else if (num==16'd16057) begin
		isPrime = 1;
	end	else if (num==16'd16061) begin
		isPrime = 1;
	end	else if (num==16'd16063) begin
		isPrime = 1;
	end	else if (num==16'd16067) begin
		isPrime = 1;
	end	else if (num==16'd16069) begin
		isPrime = 1;
	end	else if (num==16'd16073) begin
		isPrime = 1;
	end	else if (num==16'd16087) begin
		isPrime = 1;
	end	else if (num==16'd16091) begin
		isPrime = 1;
	end	else if (num==16'd16097) begin
		isPrime = 1;
	end	else if (num==16'd16103) begin
		isPrime = 1;
	end	else if (num==16'd16111) begin
		isPrime = 1;
	end	else if (num==16'd16127) begin
		isPrime = 1;
	end	else if (num==16'd16139) begin
		isPrime = 1;
	end	else if (num==16'd16141) begin
		isPrime = 1;
	end	else if (num==16'd16183) begin
		isPrime = 1;
	end	else if (num==16'd16187) begin
		isPrime = 1;
	end	else if (num==16'd16189) begin
		isPrime = 1;
	end	else if (num==16'd16193) begin
		isPrime = 1;
	end	else if (num==16'd16217) begin
		isPrime = 1;
	end	else if (num==16'd16223) begin
		isPrime = 1;
	end	else if (num==16'd16229) begin
		isPrime = 1;
	end	else if (num==16'd16231) begin
		isPrime = 1;
	end	else if (num==16'd16249) begin
		isPrime = 1;
	end	else if (num==16'd16253) begin
		isPrime = 1;
	end	else if (num==16'd16267) begin
		isPrime = 1;
	end	else if (num==16'd16273) begin
		isPrime = 1;
	end	else if (num==16'd16301) begin
		isPrime = 1;
	end	else if (num==16'd16319) begin
		isPrime = 1;
	end	else if (num==16'd16333) begin
		isPrime = 1;
	end	else if (num==16'd16339) begin
		isPrime = 1;
	end	else if (num==16'd16349) begin
		isPrime = 1;
	end	else if (num==16'd16361) begin
		isPrime = 1;
	end	else if (num==16'd16363) begin
		isPrime = 1;
	end	else if (num==16'd16369) begin
		isPrime = 1;
	end	else if (num==16'd16381) begin
		isPrime = 1;
	end	else if (num==16'd16411) begin
		isPrime = 1;
	end	else if (num==16'd16417) begin
		isPrime = 1;
	end	else if (num==16'd16421) begin
		isPrime = 1;
	end	else if (num==16'd16427) begin
		isPrime = 1;
	end	else if (num==16'd16433) begin
		isPrime = 1;
	end	else if (num==16'd16447) begin
		isPrime = 1;
	end	else if (num==16'd16451) begin
		isPrime = 1;
	end	else if (num==16'd16453) begin
		isPrime = 1;
	end	else if (num==16'd16477) begin
		isPrime = 1;
	end	else if (num==16'd16481) begin
		isPrime = 1;
	end	else if (num==16'd16487) begin
		isPrime = 1;
	end	else if (num==16'd16493) begin
		isPrime = 1;
	end	else if (num==16'd16519) begin
		isPrime = 1;
	end	else if (num==16'd16529) begin
		isPrime = 1;
	end	else if (num==16'd16547) begin
		isPrime = 1;
	end	else if (num==16'd16553) begin
		isPrime = 1;
	end	else if (num==16'd16561) begin
		isPrime = 1;
	end	else if (num==16'd16567) begin
		isPrime = 1;
	end	else if (num==16'd16573) begin
		isPrime = 1;
	end	else if (num==16'd16603) begin
		isPrime = 1;
	end	else if (num==16'd16607) begin
		isPrime = 1;
	end	else if (num==16'd16619) begin
		isPrime = 1;
	end	else if (num==16'd16631) begin
		isPrime = 1;
	end	else if (num==16'd16633) begin
		isPrime = 1;
	end	else if (num==16'd16649) begin
		isPrime = 1;
	end	else if (num==16'd16651) begin
		isPrime = 1;
	end	else if (num==16'd16657) begin
		isPrime = 1;
	end	else if (num==16'd16661) begin
		isPrime = 1;
	end	else if (num==16'd16673) begin
		isPrime = 1;
	end	else if (num==16'd16691) begin
		isPrime = 1;
	end	else if (num==16'd16693) begin
		isPrime = 1;
	end	else if (num==16'd16699) begin
		isPrime = 1;
	end	else if (num==16'd16703) begin
		isPrime = 1;
	end	else if (num==16'd16729) begin
		isPrime = 1;
	end	else if (num==16'd16741) begin
		isPrime = 1;
	end	else if (num==16'd16747) begin
		isPrime = 1;
	end	else if (num==16'd16759) begin
		isPrime = 1;
	end	else if (num==16'd16763) begin
		isPrime = 1;
	end	else if (num==16'd16787) begin
		isPrime = 1;
	end	else if (num==16'd16811) begin
		isPrime = 1;
	end	else if (num==16'd16823) begin
		isPrime = 1;
	end	else if (num==16'd16829) begin
		isPrime = 1;
	end	else if (num==16'd16831) begin
		isPrime = 1;
	end	else if (num==16'd16843) begin
		isPrime = 1;
	end	else if (num==16'd16871) begin
		isPrime = 1;
	end	else if (num==16'd16879) begin
		isPrime = 1;
	end	else if (num==16'd16883) begin
		isPrime = 1;
	end	else if (num==16'd16889) begin
		isPrime = 1;
	end	else if (num==16'd16901) begin
		isPrime = 1;
	end	else if (num==16'd16903) begin
		isPrime = 1;
	end	else if (num==16'd16921) begin
		isPrime = 1;
	end	else if (num==16'd16927) begin
		isPrime = 1;
	end	else if (num==16'd16931) begin
		isPrime = 1;
	end	else if (num==16'd16937) begin
		isPrime = 1;
	end	else if (num==16'd16943) begin
		isPrime = 1;
	end	else if (num==16'd16963) begin
		isPrime = 1;
	end	else if (num==16'd16979) begin
		isPrime = 1;
	end	else if (num==16'd16981) begin
		isPrime = 1;
	end	else if (num==16'd16987) begin
		isPrime = 1;
	end	else if (num==16'd16993) begin
		isPrime = 1;
	end	else if (num==16'd17011) begin
		isPrime = 1;
	end	else if (num==16'd17021) begin
		isPrime = 1;
	end	else if (num==16'd17027) begin
		isPrime = 1;
	end	else if (num==16'd17029) begin
		isPrime = 1;
	end	else if (num==16'd17033) begin
		isPrime = 1;
	end	else if (num==16'd17041) begin
		isPrime = 1;
	end	else if (num==16'd17047) begin
		isPrime = 1;
	end	else if (num==16'd17053) begin
		isPrime = 1;
	end	else if (num==16'd17077) begin
		isPrime = 1;
	end	else if (num==16'd17093) begin
		isPrime = 1;
	end	else if (num==16'd17099) begin
		isPrime = 1;
	end	else if (num==16'd17107) begin
		isPrime = 1;
	end	else if (num==16'd17117) begin
		isPrime = 1;
	end	else if (num==16'd17123) begin
		isPrime = 1;
	end	else if (num==16'd17137) begin
		isPrime = 1;
	end	else if (num==16'd17159) begin
		isPrime = 1;
	end	else if (num==16'd17167) begin
		isPrime = 1;
	end	else if (num==16'd17183) begin
		isPrime = 1;
	end	else if (num==16'd17189) begin
		isPrime = 1;
	end	else if (num==16'd17191) begin
		isPrime = 1;
	end	else if (num==16'd17203) begin
		isPrime = 1;
	end	else if (num==16'd17207) begin
		isPrime = 1;
	end	else if (num==16'd17209) begin
		isPrime = 1;
	end	else if (num==16'd17231) begin
		isPrime = 1;
	end	else if (num==16'd17239) begin
		isPrime = 1;
	end	else if (num==16'd17257) begin
		isPrime = 1;
	end	else if (num==16'd17291) begin
		isPrime = 1;
	end	else if (num==16'd17293) begin
		isPrime = 1;
	end	else if (num==16'd17299) begin
		isPrime = 1;
	end	else if (num==16'd17317) begin
		isPrime = 1;
	end	else if (num==16'd17321) begin
		isPrime = 1;
	end	else if (num==16'd17327) begin
		isPrime = 1;
	end	else if (num==16'd17333) begin
		isPrime = 1;
	end	else if (num==16'd17341) begin
		isPrime = 1;
	end	else if (num==16'd17351) begin
		isPrime = 1;
	end	else if (num==16'd17359) begin
		isPrime = 1;
	end	else if (num==16'd17377) begin
		isPrime = 1;
	end	else if (num==16'd17383) begin
		isPrime = 1;
	end	else if (num==16'd17387) begin
		isPrime = 1;
	end	else if (num==16'd17389) begin
		isPrime = 1;
	end	else if (num==16'd17393) begin
		isPrime = 1;
	end	else if (num==16'd17401) begin
		isPrime = 1;
	end	else if (num==16'd17417) begin
		isPrime = 1;
	end	else if (num==16'd17419) begin
		isPrime = 1;
	end	else if (num==16'd17431) begin
		isPrime = 1;
	end	else if (num==16'd17443) begin
		isPrime = 1;
	end	else if (num==16'd17449) begin
		isPrime = 1;
	end	else if (num==16'd17467) begin
		isPrime = 1;
	end	else if (num==16'd17471) begin
		isPrime = 1;
	end	else if (num==16'd17477) begin
		isPrime = 1;
	end	else if (num==16'd17483) begin
		isPrime = 1;
	end	else if (num==16'd17489) begin
		isPrime = 1;
	end	else if (num==16'd17491) begin
		isPrime = 1;
	end	else if (num==16'd17497) begin
		isPrime = 1;
	end	else if (num==16'd17509) begin
		isPrime = 1;
	end	else if (num==16'd17519) begin
		isPrime = 1;
	end	else if (num==16'd17539) begin
		isPrime = 1;
	end	else if (num==16'd17551) begin
		isPrime = 1;
	end	else if (num==16'd17569) begin
		isPrime = 1;
	end	else if (num==16'd17573) begin
		isPrime = 1;
	end	else if (num==16'd17579) begin
		isPrime = 1;
	end	else if (num==16'd17581) begin
		isPrime = 1;
	end	else if (num==16'd17597) begin
		isPrime = 1;
	end	else if (num==16'd17599) begin
		isPrime = 1;
	end	else if (num==16'd17609) begin
		isPrime = 1;
	end	else if (num==16'd17623) begin
		isPrime = 1;
	end	else if (num==16'd17627) begin
		isPrime = 1;
	end	else if (num==16'd17657) begin
		isPrime = 1;
	end	else if (num==16'd17659) begin
		isPrime = 1;
	end	else if (num==16'd17669) begin
		isPrime = 1;
	end	else if (num==16'd17681) begin
		isPrime = 1;
	end	else if (num==16'd17683) begin
		isPrime = 1;
	end	else if (num==16'd17707) begin
		isPrime = 1;
	end	else if (num==16'd17713) begin
		isPrime = 1;
	end	else if (num==16'd17729) begin
		isPrime = 1;
	end	else if (num==16'd17737) begin
		isPrime = 1;
	end	else if (num==16'd17747) begin
		isPrime = 1;
	end	else if (num==16'd17749) begin
		isPrime = 1;
	end	else if (num==16'd17761) begin
		isPrime = 1;
	end	else if (num==16'd17783) begin
		isPrime = 1;
	end	else if (num==16'd17789) begin
		isPrime = 1;
	end	else if (num==16'd17791) begin
		isPrime = 1;
	end	else if (num==16'd17807) begin
		isPrime = 1;
	end	else if (num==16'd17827) begin
		isPrime = 1;
	end	else if (num==16'd17837) begin
		isPrime = 1;
	end	else if (num==16'd17839) begin
		isPrime = 1;
	end	else if (num==16'd17851) begin
		isPrime = 1;
	end	else if (num==16'd17863) begin
		isPrime = 1;
	end	else if (num==16'd17881) begin
		isPrime = 1;
	end	else if (num==16'd17891) begin
		isPrime = 1;
	end	else if (num==16'd17903) begin
		isPrime = 1;
	end	else if (num==16'd17909) begin
		isPrime = 1;
	end	else if (num==16'd17911) begin
		isPrime = 1;
	end	else if (num==16'd17921) begin
		isPrime = 1;
	end	else if (num==16'd17923) begin
		isPrime = 1;
	end	else if (num==16'd17929) begin
		isPrime = 1;
	end	else if (num==16'd17939) begin
		isPrime = 1;
	end	else if (num==16'd17957) begin
		isPrime = 1;
	end	else if (num==16'd17959) begin
		isPrime = 1;
	end	else if (num==16'd17971) begin
		isPrime = 1;
	end	else if (num==16'd17977) begin
		isPrime = 1;
	end	else if (num==16'd17981) begin
		isPrime = 1;
	end	else if (num==16'd17987) begin
		isPrime = 1;
	end	else if (num==16'd17989) begin
		isPrime = 1;
	end	else if (num==16'd18013) begin
		isPrime = 1;
	end	else if (num==16'd18041) begin
		isPrime = 1;
	end	else if (num==16'd18043) begin
		isPrime = 1;
	end	else if (num==16'd18047) begin
		isPrime = 1;
	end	else if (num==16'd18049) begin
		isPrime = 1;
	end	else if (num==16'd18059) begin
		isPrime = 1;
	end	else if (num==16'd18061) begin
		isPrime = 1;
	end	else if (num==16'd18077) begin
		isPrime = 1;
	end	else if (num==16'd18089) begin
		isPrime = 1;
	end	else if (num==16'd18097) begin
		isPrime = 1;
	end	else if (num==16'd18119) begin
		isPrime = 1;
	end	else if (num==16'd18121) begin
		isPrime = 1;
	end	else if (num==16'd18127) begin
		isPrime = 1;
	end	else if (num==16'd18131) begin
		isPrime = 1;
	end	else if (num==16'd18133) begin
		isPrime = 1;
	end	else if (num==16'd18143) begin
		isPrime = 1;
	end	else if (num==16'd18149) begin
		isPrime = 1;
	end	else if (num==16'd18169) begin
		isPrime = 1;
	end	else if (num==16'd18181) begin
		isPrime = 1;
	end	else if (num==16'd18191) begin
		isPrime = 1;
	end	else if (num==16'd18199) begin
		isPrime = 1;
	end	else if (num==16'd18211) begin
		isPrime = 1;
	end	else if (num==16'd18217) begin
		isPrime = 1;
	end	else if (num==16'd18223) begin
		isPrime = 1;
	end	else if (num==16'd18229) begin
		isPrime = 1;
	end	else if (num==16'd18233) begin
		isPrime = 1;
	end	else if (num==16'd18251) begin
		isPrime = 1;
	end	else if (num==16'd18253) begin
		isPrime = 1;
	end	else if (num==16'd18257) begin
		isPrime = 1;
	end	else if (num==16'd18269) begin
		isPrime = 1;
	end	else if (num==16'd18287) begin
		isPrime = 1;
	end	else if (num==16'd18289) begin
		isPrime = 1;
	end	else if (num==16'd18301) begin
		isPrime = 1;
	end	else if (num==16'd18307) begin
		isPrime = 1;
	end	else if (num==16'd18311) begin
		isPrime = 1;
	end	else if (num==16'd18313) begin
		isPrime = 1;
	end	else if (num==16'd18329) begin
		isPrime = 1;
	end	else if (num==16'd18341) begin
		isPrime = 1;
	end	else if (num==16'd18353) begin
		isPrime = 1;
	end	else if (num==16'd18367) begin
		isPrime = 1;
	end	else if (num==16'd18371) begin
		isPrime = 1;
	end	else if (num==16'd18379) begin
		isPrime = 1;
	end	else if (num==16'd18397) begin
		isPrime = 1;
	end	else if (num==16'd18401) begin
		isPrime = 1;
	end	else if (num==16'd18413) begin
		isPrime = 1;
	end	else if (num==16'd18427) begin
		isPrime = 1;
	end	else if (num==16'd18433) begin
		isPrime = 1;
	end	else if (num==16'd18439) begin
		isPrime = 1;
	end	else if (num==16'd18443) begin
		isPrime = 1;
	end	else if (num==16'd18451) begin
		isPrime = 1;
	end	else if (num==16'd18457) begin
		isPrime = 1;
	end	else if (num==16'd18461) begin
		isPrime = 1;
	end	else if (num==16'd18481) begin
		isPrime = 1;
	end	else if (num==16'd18493) begin
		isPrime = 1;
	end	else if (num==16'd18503) begin
		isPrime = 1;
	end	else if (num==16'd18517) begin
		isPrime = 1;
	end	else if (num==16'd18521) begin
		isPrime = 1;
	end	else if (num==16'd18523) begin
		isPrime = 1;
	end	else if (num==16'd18539) begin
		isPrime = 1;
	end	else if (num==16'd18541) begin
		isPrime = 1;
	end	else if (num==16'd18553) begin
		isPrime = 1;
	end	else if (num==16'd18583) begin
		isPrime = 1;
	end	else if (num==16'd18587) begin
		isPrime = 1;
	end	else if (num==16'd18593) begin
		isPrime = 1;
	end	else if (num==16'd18617) begin
		isPrime = 1;
	end	else if (num==16'd18637) begin
		isPrime = 1;
	end	else if (num==16'd18661) begin
		isPrime = 1;
	end	else if (num==16'd18671) begin
		isPrime = 1;
	end	else if (num==16'd18679) begin
		isPrime = 1;
	end	else if (num==16'd18691) begin
		isPrime = 1;
	end	else if (num==16'd18701) begin
		isPrime = 1;
	end	else if (num==16'd18713) begin
		isPrime = 1;
	end	else if (num==16'd18719) begin
		isPrime = 1;
	end	else if (num==16'd18731) begin
		isPrime = 1;
	end	else if (num==16'd18743) begin
		isPrime = 1;
	end	else if (num==16'd18749) begin
		isPrime = 1;
	end	else if (num==16'd18757) begin
		isPrime = 1;
	end	else if (num==16'd18773) begin
		isPrime = 1;
	end	else if (num==16'd18787) begin
		isPrime = 1;
	end	else if (num==16'd18793) begin
		isPrime = 1;
	end	else if (num==16'd18797) begin
		isPrime = 1;
	end	else if (num==16'd18803) begin
		isPrime = 1;
	end	else if (num==16'd18839) begin
		isPrime = 1;
	end	else if (num==16'd18859) begin
		isPrime = 1;
	end	else if (num==16'd18869) begin
		isPrime = 1;
	end	else if (num==16'd18899) begin
		isPrime = 1;
	end	else if (num==16'd18911) begin
		isPrime = 1;
	end	else if (num==16'd18913) begin
		isPrime = 1;
	end	else if (num==16'd18917) begin
		isPrime = 1;
	end	else if (num==16'd18919) begin
		isPrime = 1;
	end	else if (num==16'd18947) begin
		isPrime = 1;
	end	else if (num==16'd18959) begin
		isPrime = 1;
	end	else if (num==16'd18973) begin
		isPrime = 1;
	end	else if (num==16'd18979) begin
		isPrime = 1;
	end	else if (num==16'd19001) begin
		isPrime = 1;
	end	else if (num==16'd19009) begin
		isPrime = 1;
	end	else if (num==16'd19013) begin
		isPrime = 1;
	end	else if (num==16'd19031) begin
		isPrime = 1;
	end	else if (num==16'd19037) begin
		isPrime = 1;
	end	else if (num==16'd19051) begin
		isPrime = 1;
	end	else if (num==16'd19069) begin
		isPrime = 1;
	end	else if (num==16'd19073) begin
		isPrime = 1;
	end	else if (num==16'd19079) begin
		isPrime = 1;
	end	else if (num==16'd19081) begin
		isPrime = 1;
	end	else if (num==16'd19087) begin
		isPrime = 1;
	end	else if (num==16'd19121) begin
		isPrime = 1;
	end	else if (num==16'd19139) begin
		isPrime = 1;
	end	else if (num==16'd19141) begin
		isPrime = 1;
	end	else if (num==16'd19157) begin
		isPrime = 1;
	end	else if (num==16'd19163) begin
		isPrime = 1;
	end	else if (num==16'd19181) begin
		isPrime = 1;
	end	else if (num==16'd19183) begin
		isPrime = 1;
	end	else if (num==16'd19207) begin
		isPrime = 1;
	end	else if (num==16'd19211) begin
		isPrime = 1;
	end	else if (num==16'd19213) begin
		isPrime = 1;
	end	else if (num==16'd19219) begin
		isPrime = 1;
	end	else if (num==16'd19231) begin
		isPrime = 1;
	end	else if (num==16'd19237) begin
		isPrime = 1;
	end	else if (num==16'd19249) begin
		isPrime = 1;
	end	else if (num==16'd19259) begin
		isPrime = 1;
	end	else if (num==16'd19267) begin
		isPrime = 1;
	end	else if (num==16'd19273) begin
		isPrime = 1;
	end	else if (num==16'd19289) begin
		isPrime = 1;
	end	else if (num==16'd19301) begin
		isPrime = 1;
	end	else if (num==16'd19309) begin
		isPrime = 1;
	end	else if (num==16'd19319) begin
		isPrime = 1;
	end	else if (num==16'd19333) begin
		isPrime = 1;
	end	else if (num==16'd19373) begin
		isPrime = 1;
	end	else if (num==16'd19379) begin
		isPrime = 1;
	end	else if (num==16'd19381) begin
		isPrime = 1;
	end	else if (num==16'd19387) begin
		isPrime = 1;
	end	else if (num==16'd19391) begin
		isPrime = 1;
	end	else if (num==16'd19403) begin
		isPrime = 1;
	end	else if (num==16'd19417) begin
		isPrime = 1;
	end	else if (num==16'd19421) begin
		isPrime = 1;
	end	else if (num==16'd19423) begin
		isPrime = 1;
	end	else if (num==16'd19427) begin
		isPrime = 1;
	end	else if (num==16'd19429) begin
		isPrime = 1;
	end	else if (num==16'd19433) begin
		isPrime = 1;
	end	else if (num==16'd19441) begin
		isPrime = 1;
	end	else if (num==16'd19447) begin
		isPrime = 1;
	end	else if (num==16'd19457) begin
		isPrime = 1;
	end	else if (num==16'd19463) begin
		isPrime = 1;
	end	else if (num==16'd19469) begin
		isPrime = 1;
	end	else if (num==16'd19471) begin
		isPrime = 1;
	end	else if (num==16'd19477) begin
		isPrime = 1;
	end	else if (num==16'd19483) begin
		isPrime = 1;
	end	else if (num==16'd19489) begin
		isPrime = 1;
	end	else if (num==16'd19501) begin
		isPrime = 1;
	end	else if (num==16'd19507) begin
		isPrime = 1;
	end	else if (num==16'd19531) begin
		isPrime = 1;
	end	else if (num==16'd19541) begin
		isPrime = 1;
	end	else if (num==16'd19543) begin
		isPrime = 1;
	end	else if (num==16'd19553) begin
		isPrime = 1;
	end	else if (num==16'd19559) begin
		isPrime = 1;
	end	else if (num==16'd19571) begin
		isPrime = 1;
	end	else if (num==16'd19577) begin
		isPrime = 1;
	end	else if (num==16'd19583) begin
		isPrime = 1;
	end	else if (num==16'd19597) begin
		isPrime = 1;
	end	else if (num==16'd19603) begin
		isPrime = 1;
	end	else if (num==16'd19609) begin
		isPrime = 1;
	end	else if (num==16'd19661) begin
		isPrime = 1;
	end	else if (num==16'd19681) begin
		isPrime = 1;
	end	else if (num==16'd19687) begin
		isPrime = 1;
	end	else if (num==16'd19697) begin
		isPrime = 1;
	end	else if (num==16'd19699) begin
		isPrime = 1;
	end	else if (num==16'd19709) begin
		isPrime = 1;
	end	else if (num==16'd19717) begin
		isPrime = 1;
	end	else if (num==16'd19727) begin
		isPrime = 1;
	end	else if (num==16'd19739) begin
		isPrime = 1;
	end	else if (num==16'd19751) begin
		isPrime = 1;
	end	else if (num==16'd19753) begin
		isPrime = 1;
	end	else if (num==16'd19759) begin
		isPrime = 1;
	end	else if (num==16'd19763) begin
		isPrime = 1;
	end	else if (num==16'd19777) begin
		isPrime = 1;
	end	else if (num==16'd19793) begin
		isPrime = 1;
	end	else if (num==16'd19801) begin
		isPrime = 1;
	end	else if (num==16'd19813) begin
		isPrime = 1;
	end	else if (num==16'd19819) begin
		isPrime = 1;
	end	else if (num==16'd19841) begin
		isPrime = 1;
	end	else if (num==16'd19843) begin
		isPrime = 1;
	end	else if (num==16'd19853) begin
		isPrime = 1;
	end	else if (num==16'd19861) begin
		isPrime = 1;
	end	else if (num==16'd19867) begin
		isPrime = 1;
	end	else if (num==16'd19889) begin
		isPrime = 1;
	end	else if (num==16'd19891) begin
		isPrime = 1;
	end	else if (num==16'd19913) begin
		isPrime = 1;
	end	else if (num==16'd19919) begin
		isPrime = 1;
	end	else if (num==16'd19927) begin
		isPrime = 1;
	end	else if (num==16'd19937) begin
		isPrime = 1;
	end	else if (num==16'd19949) begin
		isPrime = 1;
	end	else if (num==16'd19961) begin
		isPrime = 1;
	end	else if (num==16'd19963) begin
		isPrime = 1;
	end	else if (num==16'd19973) begin
		isPrime = 1;
	end	else if (num==16'd19979) begin
		isPrime = 1;
	end	else if (num==16'd19991) begin
		isPrime = 1;
	end	else if (num==16'd19993) begin
		isPrime = 1;
	end	else if (num==16'd19997) begin
		isPrime = 1;
	end	else if (num==16'd20011) begin
		isPrime = 1;
	end	else if (num==16'd20021) begin
		isPrime = 1;
	end	else if (num==16'd20023) begin
		isPrime = 1;
	end	else if (num==16'd20029) begin
		isPrime = 1;
	end	else if (num==16'd20047) begin
		isPrime = 1;
	end	else if (num==16'd20051) begin
		isPrime = 1;
	end	else if (num==16'd20063) begin
		isPrime = 1;
	end	else if (num==16'd20071) begin
		isPrime = 1;
	end	else if (num==16'd20089) begin
		isPrime = 1;
	end	else if (num==16'd20101) begin
		isPrime = 1;
	end	else if (num==16'd20107) begin
		isPrime = 1;
	end	else if (num==16'd20113) begin
		isPrime = 1;
	end	else if (num==16'd20117) begin
		isPrime = 1;
	end	else if (num==16'd20123) begin
		isPrime = 1;
	end	else if (num==16'd20129) begin
		isPrime = 1;
	end	else if (num==16'd20143) begin
		isPrime = 1;
	end	else if (num==16'd20147) begin
		isPrime = 1;
	end	else if (num==16'd20149) begin
		isPrime = 1;
	end	else if (num==16'd20161) begin
		isPrime = 1;
	end	else if (num==16'd20173) begin
		isPrime = 1;
	end	else if (num==16'd20177) begin
		isPrime = 1;
	end	else if (num==16'd20183) begin
		isPrime = 1;
	end	else if (num==16'd20201) begin
		isPrime = 1;
	end	else if (num==16'd20219) begin
		isPrime = 1;
	end	else if (num==16'd20231) begin
		isPrime = 1;
	end	else if (num==16'd20233) begin
		isPrime = 1;
	end	else if (num==16'd20249) begin
		isPrime = 1;
	end	else if (num==16'd20261) begin
		isPrime = 1;
	end	else if (num==16'd20269) begin
		isPrime = 1;
	end	else if (num==16'd20287) begin
		isPrime = 1;
	end	else if (num==16'd20297) begin
		isPrime = 1;
	end	else if (num==16'd20323) begin
		isPrime = 1;
	end	else if (num==16'd20327) begin
		isPrime = 1;
	end	else if (num==16'd20333) begin
		isPrime = 1;
	end	else if (num==16'd20341) begin
		isPrime = 1;
	end	else if (num==16'd20347) begin
		isPrime = 1;
	end	else if (num==16'd20353) begin
		isPrime = 1;
	end	else if (num==16'd20357) begin
		isPrime = 1;
	end	else if (num==16'd20359) begin
		isPrime = 1;
	end	else if (num==16'd20369) begin
		isPrime = 1;
	end	else if (num==16'd20389) begin
		isPrime = 1;
	end	else if (num==16'd20393) begin
		isPrime = 1;
	end	else if (num==16'd20399) begin
		isPrime = 1;
	end	else if (num==16'd20407) begin
		isPrime = 1;
	end	else if (num==16'd20411) begin
		isPrime = 1;
	end	else if (num==16'd20431) begin
		isPrime = 1;
	end	else if (num==16'd20441) begin
		isPrime = 1;
	end	else if (num==16'd20443) begin
		isPrime = 1;
	end	else if (num==16'd20477) begin
		isPrime = 1;
	end	else if (num==16'd20479) begin
		isPrime = 1;
	end	else if (num==16'd20483) begin
		isPrime = 1;
	end	else if (num==16'd20507) begin
		isPrime = 1;
	end	else if (num==16'd20509) begin
		isPrime = 1;
	end	else if (num==16'd20521) begin
		isPrime = 1;
	end	else if (num==16'd20533) begin
		isPrime = 1;
	end	else if (num==16'd20543) begin
		isPrime = 1;
	end	else if (num==16'd20549) begin
		isPrime = 1;
	end	else if (num==16'd20551) begin
		isPrime = 1;
	end	else if (num==16'd20563) begin
		isPrime = 1;
	end	else if (num==16'd20593) begin
		isPrime = 1;
	end	else if (num==16'd20599) begin
		isPrime = 1;
	end	else if (num==16'd20611) begin
		isPrime = 1;
	end	else if (num==16'd20627) begin
		isPrime = 1;
	end	else if (num==16'd20639) begin
		isPrime = 1;
	end	else if (num==16'd20641) begin
		isPrime = 1;
	end	else if (num==16'd20663) begin
		isPrime = 1;
	end	else if (num==16'd20681) begin
		isPrime = 1;
	end	else if (num==16'd20693) begin
		isPrime = 1;
	end	else if (num==16'd20707) begin
		isPrime = 1;
	end	else if (num==16'd20717) begin
		isPrime = 1;
	end	else if (num==16'd20719) begin
		isPrime = 1;
	end	else if (num==16'd20731) begin
		isPrime = 1;
	end	else if (num==16'd20743) begin
		isPrime = 1;
	end	else if (num==16'd20747) begin
		isPrime = 1;
	end	else if (num==16'd20749) begin
		isPrime = 1;
	end	else if (num==16'd20753) begin
		isPrime = 1;
	end	else if (num==16'd20759) begin
		isPrime = 1;
	end	else if (num==16'd20771) begin
		isPrime = 1;
	end	else if (num==16'd20773) begin
		isPrime = 1;
	end	else if (num==16'd20789) begin
		isPrime = 1;
	end	else if (num==16'd20807) begin
		isPrime = 1;
	end	else if (num==16'd20809) begin
		isPrime = 1;
	end	else if (num==16'd20849) begin
		isPrime = 1;
	end	else if (num==16'd20857) begin
		isPrime = 1;
	end	else if (num==16'd20873) begin
		isPrime = 1;
	end	else if (num==16'd20879) begin
		isPrime = 1;
	end	else if (num==16'd20887) begin
		isPrime = 1;
	end	else if (num==16'd20897) begin
		isPrime = 1;
	end	else if (num==16'd20899) begin
		isPrime = 1;
	end	else if (num==16'd20903) begin
		isPrime = 1;
	end	else if (num==16'd20921) begin
		isPrime = 1;
	end	else if (num==16'd20929) begin
		isPrime = 1;
	end	else if (num==16'd20939) begin
		isPrime = 1;
	end	else if (num==16'd20947) begin
		isPrime = 1;
	end	else if (num==16'd20959) begin
		isPrime = 1;
	end	else if (num==16'd20963) begin
		isPrime = 1;
	end	else if (num==16'd20981) begin
		isPrime = 1;
	end	else if (num==16'd20983) begin
		isPrime = 1;
	end	else if (num==16'd21001) begin
		isPrime = 1;
	end	else if (num==16'd21011) begin
		isPrime = 1;
	end	else if (num==16'd21013) begin
		isPrime = 1;
	end	else if (num==16'd21017) begin
		isPrime = 1;
	end	else if (num==16'd21019) begin
		isPrime = 1;
	end	else if (num==16'd21023) begin
		isPrime = 1;
	end	else if (num==16'd21031) begin
		isPrime = 1;
	end	else if (num==16'd21059) begin
		isPrime = 1;
	end	else if (num==16'd21061) begin
		isPrime = 1;
	end	else if (num==16'd21067) begin
		isPrime = 1;
	end	else if (num==16'd21089) begin
		isPrime = 1;
	end	else if (num==16'd21101) begin
		isPrime = 1;
	end	else if (num==16'd21107) begin
		isPrime = 1;
	end	else if (num==16'd21121) begin
		isPrime = 1;
	end	else if (num==16'd21139) begin
		isPrime = 1;
	end	else if (num==16'd21143) begin
		isPrime = 1;
	end	else if (num==16'd21149) begin
		isPrime = 1;
	end	else if (num==16'd21157) begin
		isPrime = 1;
	end	else if (num==16'd21163) begin
		isPrime = 1;
	end	else if (num==16'd21169) begin
		isPrime = 1;
	end	else if (num==16'd21179) begin
		isPrime = 1;
	end	else if (num==16'd21187) begin
		isPrime = 1;
	end	else if (num==16'd21191) begin
		isPrime = 1;
	end	else if (num==16'd21193) begin
		isPrime = 1;
	end	else if (num==16'd21211) begin
		isPrime = 1;
	end	else if (num==16'd21221) begin
		isPrime = 1;
	end	else if (num==16'd21227) begin
		isPrime = 1;
	end	else if (num==16'd21247) begin
		isPrime = 1;
	end	else if (num==16'd21269) begin
		isPrime = 1;
	end	else if (num==16'd21277) begin
		isPrime = 1;
	end	else if (num==16'd21283) begin
		isPrime = 1;
	end	else if (num==16'd21313) begin
		isPrime = 1;
	end	else if (num==16'd21317) begin
		isPrime = 1;
	end	else if (num==16'd21319) begin
		isPrime = 1;
	end	else if (num==16'd21323) begin
		isPrime = 1;
	end	else if (num==16'd21341) begin
		isPrime = 1;
	end	else if (num==16'd21347) begin
		isPrime = 1;
	end	else if (num==16'd21377) begin
		isPrime = 1;
	end	else if (num==16'd21379) begin
		isPrime = 1;
	end	else if (num==16'd21383) begin
		isPrime = 1;
	end	else if (num==16'd21391) begin
		isPrime = 1;
	end	else if (num==16'd21397) begin
		isPrime = 1;
	end	else if (num==16'd21401) begin
		isPrime = 1;
	end	else if (num==16'd21407) begin
		isPrime = 1;
	end	else if (num==16'd21419) begin
		isPrime = 1;
	end	else if (num==16'd21433) begin
		isPrime = 1;
	end	else if (num==16'd21467) begin
		isPrime = 1;
	end	else if (num==16'd21481) begin
		isPrime = 1;
	end	else if (num==16'd21487) begin
		isPrime = 1;
	end	else if (num==16'd21491) begin
		isPrime = 1;
	end	else if (num==16'd21493) begin
		isPrime = 1;
	end	else if (num==16'd21499) begin
		isPrime = 1;
	end	else if (num==16'd21503) begin
		isPrime = 1;
	end	else if (num==16'd21517) begin
		isPrime = 1;
	end	else if (num==16'd21521) begin
		isPrime = 1;
	end	else if (num==16'd21523) begin
		isPrime = 1;
	end	else if (num==16'd21529) begin
		isPrime = 1;
	end	else if (num==16'd21557) begin
		isPrime = 1;
	end	else if (num==16'd21559) begin
		isPrime = 1;
	end	else if (num==16'd21563) begin
		isPrime = 1;
	end	else if (num==16'd21569) begin
		isPrime = 1;
	end	else if (num==16'd21577) begin
		isPrime = 1;
	end	else if (num==16'd21587) begin
		isPrime = 1;
	end	else if (num==16'd21589) begin
		isPrime = 1;
	end	else if (num==16'd21599) begin
		isPrime = 1;
	end	else if (num==16'd21601) begin
		isPrime = 1;
	end	else if (num==16'd21611) begin
		isPrime = 1;
	end	else if (num==16'd21613) begin
		isPrime = 1;
	end	else if (num==16'd21617) begin
		isPrime = 1;
	end	else if (num==16'd21647) begin
		isPrime = 1;
	end	else if (num==16'd21649) begin
		isPrime = 1;
	end	else if (num==16'd21661) begin
		isPrime = 1;
	end	else if (num==16'd21673) begin
		isPrime = 1;
	end	else if (num==16'd21683) begin
		isPrime = 1;
	end	else if (num==16'd21701) begin
		isPrime = 1;
	end	else if (num==16'd21713) begin
		isPrime = 1;
	end	else if (num==16'd21727) begin
		isPrime = 1;
	end	else if (num==16'd21737) begin
		isPrime = 1;
	end	else if (num==16'd21739) begin
		isPrime = 1;
	end	else if (num==16'd21751) begin
		isPrime = 1;
	end	else if (num==16'd21757) begin
		isPrime = 1;
	end	else if (num==16'd21767) begin
		isPrime = 1;
	end	else if (num==16'd21773) begin
		isPrime = 1;
	end	else if (num==16'd21787) begin
		isPrime = 1;
	end	else if (num==16'd21799) begin
		isPrime = 1;
	end	else if (num==16'd21803) begin
		isPrime = 1;
	end	else if (num==16'd21817) begin
		isPrime = 1;
	end	else if (num==16'd21821) begin
		isPrime = 1;
	end	else if (num==16'd21839) begin
		isPrime = 1;
	end	else if (num==16'd21841) begin
		isPrime = 1;
	end	else if (num==16'd21851) begin
		isPrime = 1;
	end	else if (num==16'd21859) begin
		isPrime = 1;
	end	else if (num==16'd21863) begin
		isPrime = 1;
	end	else if (num==16'd21871) begin
		isPrime = 1;
	end	else if (num==16'd21881) begin
		isPrime = 1;
	end	else if (num==16'd21893) begin
		isPrime = 1;
	end	else if (num==16'd21911) begin
		isPrime = 1;
	end	else if (num==16'd21929) begin
		isPrime = 1;
	end	else if (num==16'd21937) begin
		isPrime = 1;
	end	else if (num==16'd21943) begin
		isPrime = 1;
	end	else if (num==16'd21961) begin
		isPrime = 1;
	end	else if (num==16'd21977) begin
		isPrime = 1;
	end	else if (num==16'd21991) begin
		isPrime = 1;
	end	else if (num==16'd21997) begin
		isPrime = 1;
	end	else if (num==16'd22003) begin
		isPrime = 1;
	end	else if (num==16'd22013) begin
		isPrime = 1;
	end	else if (num==16'd22027) begin
		isPrime = 1;
	end	else if (num==16'd22031) begin
		isPrime = 1;
	end	else if (num==16'd22037) begin
		isPrime = 1;
	end	else if (num==16'd22039) begin
		isPrime = 1;
	end	else if (num==16'd22051) begin
		isPrime = 1;
	end	else if (num==16'd22063) begin
		isPrime = 1;
	end	else if (num==16'd22067) begin
		isPrime = 1;
	end	else if (num==16'd22073) begin
		isPrime = 1;
	end	else if (num==16'd22079) begin
		isPrime = 1;
	end	else if (num==16'd22091) begin
		isPrime = 1;
	end	else if (num==16'd22093) begin
		isPrime = 1;
	end	else if (num==16'd22109) begin
		isPrime = 1;
	end	else if (num==16'd22111) begin
		isPrime = 1;
	end	else if (num==16'd22123) begin
		isPrime = 1;
	end	else if (num==16'd22129) begin
		isPrime = 1;
	end	else if (num==16'd22133) begin
		isPrime = 1;
	end	else if (num==16'd22147) begin
		isPrime = 1;
	end	else if (num==16'd22153) begin
		isPrime = 1;
	end	else if (num==16'd22157) begin
		isPrime = 1;
	end	else if (num==16'd22159) begin
		isPrime = 1;
	end	else if (num==16'd22171) begin
		isPrime = 1;
	end	else if (num==16'd22189) begin
		isPrime = 1;
	end	else if (num==16'd22193) begin
		isPrime = 1;
	end	else if (num==16'd22229) begin
		isPrime = 1;
	end	else if (num==16'd22247) begin
		isPrime = 1;
	end	else if (num==16'd22259) begin
		isPrime = 1;
	end	else if (num==16'd22271) begin
		isPrime = 1;
	end	else if (num==16'd22273) begin
		isPrime = 1;
	end	else if (num==16'd22277) begin
		isPrime = 1;
	end	else if (num==16'd22279) begin
		isPrime = 1;
	end	else if (num==16'd22283) begin
		isPrime = 1;
	end	else if (num==16'd22291) begin
		isPrime = 1;
	end	else if (num==16'd22303) begin
		isPrime = 1;
	end	else if (num==16'd22307) begin
		isPrime = 1;
	end	else if (num==16'd22343) begin
		isPrime = 1;
	end	else if (num==16'd22349) begin
		isPrime = 1;
	end	else if (num==16'd22367) begin
		isPrime = 1;
	end	else if (num==16'd22369) begin
		isPrime = 1;
	end	else if (num==16'd22381) begin
		isPrime = 1;
	end	else if (num==16'd22391) begin
		isPrime = 1;
	end	else if (num==16'd22397) begin
		isPrime = 1;
	end	else if (num==16'd22409) begin
		isPrime = 1;
	end	else if (num==16'd22433) begin
		isPrime = 1;
	end	else if (num==16'd22441) begin
		isPrime = 1;
	end	else if (num==16'd22447) begin
		isPrime = 1;
	end	else if (num==16'd22453) begin
		isPrime = 1;
	end	else if (num==16'd22469) begin
		isPrime = 1;
	end	else if (num==16'd22481) begin
		isPrime = 1;
	end	else if (num==16'd22483) begin
		isPrime = 1;
	end	else if (num==16'd22501) begin
		isPrime = 1;
	end	else if (num==16'd22511) begin
		isPrime = 1;
	end	else if (num==16'd22531) begin
		isPrime = 1;
	end	else if (num==16'd22541) begin
		isPrime = 1;
	end	else if (num==16'd22543) begin
		isPrime = 1;
	end	else if (num==16'd22549) begin
		isPrime = 1;
	end	else if (num==16'd22567) begin
		isPrime = 1;
	end	else if (num==16'd22571) begin
		isPrime = 1;
	end	else if (num==16'd22573) begin
		isPrime = 1;
	end	else if (num==16'd22613) begin
		isPrime = 1;
	end	else if (num==16'd22619) begin
		isPrime = 1;
	end	else if (num==16'd22621) begin
		isPrime = 1;
	end	else if (num==16'd22637) begin
		isPrime = 1;
	end	else if (num==16'd22639) begin
		isPrime = 1;
	end	else if (num==16'd22643) begin
		isPrime = 1;
	end	else if (num==16'd22651) begin
		isPrime = 1;
	end	else if (num==16'd22669) begin
		isPrime = 1;
	end	else if (num==16'd22679) begin
		isPrime = 1;
	end	else if (num==16'd22691) begin
		isPrime = 1;
	end	else if (num==16'd22697) begin
		isPrime = 1;
	end	else if (num==16'd22699) begin
		isPrime = 1;
	end	else if (num==16'd22709) begin
		isPrime = 1;
	end	else if (num==16'd22717) begin
		isPrime = 1;
	end	else if (num==16'd22721) begin
		isPrime = 1;
	end	else if (num==16'd22727) begin
		isPrime = 1;
	end	else if (num==16'd22739) begin
		isPrime = 1;
	end	else if (num==16'd22741) begin
		isPrime = 1;
	end	else if (num==16'd22751) begin
		isPrime = 1;
	end	else if (num==16'd22769) begin
		isPrime = 1;
	end	else if (num==16'd22777) begin
		isPrime = 1;
	end	else if (num==16'd22783) begin
		isPrime = 1;
	end	else if (num==16'd22787) begin
		isPrime = 1;
	end	else if (num==16'd22807) begin
		isPrime = 1;
	end	else if (num==16'd22811) begin
		isPrime = 1;
	end	else if (num==16'd22817) begin
		isPrime = 1;
	end	else if (num==16'd22853) begin
		isPrime = 1;
	end	else if (num==16'd22859) begin
		isPrime = 1;
	end	else if (num==16'd22861) begin
		isPrime = 1;
	end	else if (num==16'd22871) begin
		isPrime = 1;
	end	else if (num==16'd22877) begin
		isPrime = 1;
	end	else if (num==16'd22901) begin
		isPrime = 1;
	end	else if (num==16'd22907) begin
		isPrime = 1;
	end	else if (num==16'd22921) begin
		isPrime = 1;
	end	else if (num==16'd22937) begin
		isPrime = 1;
	end	else if (num==16'd22943) begin
		isPrime = 1;
	end	else if (num==16'd22961) begin
		isPrime = 1;
	end	else if (num==16'd22963) begin
		isPrime = 1;
	end	else if (num==16'd22973) begin
		isPrime = 1;
	end	else if (num==16'd22993) begin
		isPrime = 1;
	end	else if (num==16'd23003) begin
		isPrime = 1;
	end	else if (num==16'd23011) begin
		isPrime = 1;
	end	else if (num==16'd23017) begin
		isPrime = 1;
	end	else if (num==16'd23021) begin
		isPrime = 1;
	end	else if (num==16'd23027) begin
		isPrime = 1;
	end	else if (num==16'd23029) begin
		isPrime = 1;
	end	else if (num==16'd23039) begin
		isPrime = 1;
	end	else if (num==16'd23041) begin
		isPrime = 1;
	end	else if (num==16'd23053) begin
		isPrime = 1;
	end	else if (num==16'd23057) begin
		isPrime = 1;
	end	else if (num==16'd23059) begin
		isPrime = 1;
	end	else if (num==16'd23063) begin
		isPrime = 1;
	end	else if (num==16'd23071) begin
		isPrime = 1;
	end	else if (num==16'd23081) begin
		isPrime = 1;
	end	else if (num==16'd23087) begin
		isPrime = 1;
	end	else if (num==16'd23099) begin
		isPrime = 1;
	end	else if (num==16'd23117) begin
		isPrime = 1;
	end	else if (num==16'd23131) begin
		isPrime = 1;
	end	else if (num==16'd23143) begin
		isPrime = 1;
	end	else if (num==16'd23159) begin
		isPrime = 1;
	end	else if (num==16'd23167) begin
		isPrime = 1;
	end	else if (num==16'd23173) begin
		isPrime = 1;
	end	else if (num==16'd23189) begin
		isPrime = 1;
	end	else if (num==16'd23197) begin
		isPrime = 1;
	end	else if (num==16'd23201) begin
		isPrime = 1;
	end	else if (num==16'd23203) begin
		isPrime = 1;
	end	else if (num==16'd23209) begin
		isPrime = 1;
	end	else if (num==16'd23227) begin
		isPrime = 1;
	end	else if (num==16'd23251) begin
		isPrime = 1;
	end	else if (num==16'd23269) begin
		isPrime = 1;
	end	else if (num==16'd23279) begin
		isPrime = 1;
	end	else if (num==16'd23291) begin
		isPrime = 1;
	end	else if (num==16'd23293) begin
		isPrime = 1;
	end	else if (num==16'd23297) begin
		isPrime = 1;
	end	else if (num==16'd23311) begin
		isPrime = 1;
	end	else if (num==16'd23321) begin
		isPrime = 1;
	end	else if (num==16'd23327) begin
		isPrime = 1;
	end	else if (num==16'd23333) begin
		isPrime = 1;
	end	else if (num==16'd23339) begin
		isPrime = 1;
	end	else if (num==16'd23357) begin
		isPrime = 1;
	end	else if (num==16'd23369) begin
		isPrime = 1;
	end	else if (num==16'd23371) begin
		isPrime = 1;
	end	else if (num==16'd23399) begin
		isPrime = 1;
	end	else if (num==16'd23417) begin
		isPrime = 1;
	end	else if (num==16'd23431) begin
		isPrime = 1;
	end	else if (num==16'd23447) begin
		isPrime = 1;
	end	else if (num==16'd23459) begin
		isPrime = 1;
	end	else if (num==16'd23473) begin
		isPrime = 1;
	end	else if (num==16'd23497) begin
		isPrime = 1;
	end	else if (num==16'd23509) begin
		isPrime = 1;
	end	else if (num==16'd23531) begin
		isPrime = 1;
	end	else if (num==16'd23537) begin
		isPrime = 1;
	end	else if (num==16'd23539) begin
		isPrime = 1;
	end	else if (num==16'd23549) begin
		isPrime = 1;
	end	else if (num==16'd23557) begin
		isPrime = 1;
	end	else if (num==16'd23561) begin
		isPrime = 1;
	end	else if (num==16'd23563) begin
		isPrime = 1;
	end	else if (num==16'd23567) begin
		isPrime = 1;
	end	else if (num==16'd23581) begin
		isPrime = 1;
	end	else if (num==16'd23593) begin
		isPrime = 1;
	end	else if (num==16'd23599) begin
		isPrime = 1;
	end	else if (num==16'd23603) begin
		isPrime = 1;
	end	else if (num==16'd23609) begin
		isPrime = 1;
	end	else if (num==16'd23623) begin
		isPrime = 1;
	end	else if (num==16'd23627) begin
		isPrime = 1;
	end	else if (num==16'd23629) begin
		isPrime = 1;
	end	else if (num==16'd23633) begin
		isPrime = 1;
	end	else if (num==16'd23663) begin
		isPrime = 1;
	end	else if (num==16'd23669) begin
		isPrime = 1;
	end	else if (num==16'd23671) begin
		isPrime = 1;
	end	else if (num==16'd23677) begin
		isPrime = 1;
	end	else if (num==16'd23687) begin
		isPrime = 1;
	end	else if (num==16'd23689) begin
		isPrime = 1;
	end	else if (num==16'd23719) begin
		isPrime = 1;
	end	else if (num==16'd23741) begin
		isPrime = 1;
	end	else if (num==16'd23743) begin
		isPrime = 1;
	end	else if (num==16'd23747) begin
		isPrime = 1;
	end	else if (num==16'd23753) begin
		isPrime = 1;
	end	else if (num==16'd23761) begin
		isPrime = 1;
	end	else if (num==16'd23767) begin
		isPrime = 1;
	end	else if (num==16'd23773) begin
		isPrime = 1;
	end	else if (num==16'd23789) begin
		isPrime = 1;
	end	else if (num==16'd23801) begin
		isPrime = 1;
	end	else if (num==16'd23813) begin
		isPrime = 1;
	end	else if (num==16'd23819) begin
		isPrime = 1;
	end	else if (num==16'd23827) begin
		isPrime = 1;
	end	else if (num==16'd23831) begin
		isPrime = 1;
	end	else if (num==16'd23833) begin
		isPrime = 1;
	end	else if (num==16'd23857) begin
		isPrime = 1;
	end	else if (num==16'd23869) begin
		isPrime = 1;
	end	else if (num==16'd23873) begin
		isPrime = 1;
	end	else if (num==16'd23879) begin
		isPrime = 1;
	end	else if (num==16'd23887) begin
		isPrime = 1;
	end	else if (num==16'd23893) begin
		isPrime = 1;
	end	else if (num==16'd23899) begin
		isPrime = 1;
	end	else if (num==16'd23909) begin
		isPrime = 1;
	end	else if (num==16'd23911) begin
		isPrime = 1;
	end	else if (num==16'd23917) begin
		isPrime = 1;
	end	else if (num==16'd23929) begin
		isPrime = 1;
	end	else if (num==16'd23957) begin
		isPrime = 1;
	end	else if (num==16'd23971) begin
		isPrime = 1;
	end	else if (num==16'd23977) begin
		isPrime = 1;
	end	else if (num==16'd23981) begin
		isPrime = 1;
	end	else if (num==16'd23993) begin
		isPrime = 1;
	end	else if (num==16'd24001) begin
		isPrime = 1;
	end	else if (num==16'd24007) begin
		isPrime = 1;
	end	else if (num==16'd24019) begin
		isPrime = 1;
	end	else if (num==16'd24023) begin
		isPrime = 1;
	end	else if (num==16'd24029) begin
		isPrime = 1;
	end	else if (num==16'd24043) begin
		isPrime = 1;
	end	else if (num==16'd24049) begin
		isPrime = 1;
	end	else if (num==16'd24061) begin
		isPrime = 1;
	end	else if (num==16'd24071) begin
		isPrime = 1;
	end	else if (num==16'd24077) begin
		isPrime = 1;
	end	else if (num==16'd24083) begin
		isPrime = 1;
	end	else if (num==16'd24091) begin
		isPrime = 1;
	end	else if (num==16'd24097) begin
		isPrime = 1;
	end	else if (num==16'd24103) begin
		isPrime = 1;
	end	else if (num==16'd24107) begin
		isPrime = 1;
	end	else if (num==16'd24109) begin
		isPrime = 1;
	end	else if (num==16'd24113) begin
		isPrime = 1;
	end	else if (num==16'd24121) begin
		isPrime = 1;
	end	else if (num==16'd24133) begin
		isPrime = 1;
	end	else if (num==16'd24137) begin
		isPrime = 1;
	end	else if (num==16'd24151) begin
		isPrime = 1;
	end	else if (num==16'd24169) begin
		isPrime = 1;
	end	else if (num==16'd24179) begin
		isPrime = 1;
	end	else if (num==16'd24181) begin
		isPrime = 1;
	end	else if (num==16'd24197) begin
		isPrime = 1;
	end	else if (num==16'd24203) begin
		isPrime = 1;
	end	else if (num==16'd24223) begin
		isPrime = 1;
	end	else if (num==16'd24229) begin
		isPrime = 1;
	end	else if (num==16'd24239) begin
		isPrime = 1;
	end	else if (num==16'd24247) begin
		isPrime = 1;
	end	else if (num==16'd24251) begin
		isPrime = 1;
	end	else if (num==16'd24281) begin
		isPrime = 1;
	end	else if (num==16'd24317) begin
		isPrime = 1;
	end	else if (num==16'd24329) begin
		isPrime = 1;
	end	else if (num==16'd24337) begin
		isPrime = 1;
	end	else if (num==16'd24359) begin
		isPrime = 1;
	end	else if (num==16'd24371) begin
		isPrime = 1;
	end	else if (num==16'd24373) begin
		isPrime = 1;
	end	else if (num==16'd24379) begin
		isPrime = 1;
	end	else if (num==16'd24391) begin
		isPrime = 1;
	end	else if (num==16'd24407) begin
		isPrime = 1;
	end	else if (num==16'd24413) begin
		isPrime = 1;
	end	else if (num==16'd24419) begin
		isPrime = 1;
	end	else if (num==16'd24421) begin
		isPrime = 1;
	end	else if (num==16'd24439) begin
		isPrime = 1;
	end	else if (num==16'd24443) begin
		isPrime = 1;
	end	else if (num==16'd24469) begin
		isPrime = 1;
	end	else if (num==16'd24473) begin
		isPrime = 1;
	end	else if (num==16'd24481) begin
		isPrime = 1;
	end	else if (num==16'd24499) begin
		isPrime = 1;
	end	else if (num==16'd24509) begin
		isPrime = 1;
	end	else if (num==16'd24517) begin
		isPrime = 1;
	end	else if (num==16'd24527) begin
		isPrime = 1;
	end	else if (num==16'd24533) begin
		isPrime = 1;
	end	else if (num==16'd24547) begin
		isPrime = 1;
	end	else if (num==16'd24551) begin
		isPrime = 1;
	end	else if (num==16'd24571) begin
		isPrime = 1;
	end	else if (num==16'd24593) begin
		isPrime = 1;
	end	else if (num==16'd24611) begin
		isPrime = 1;
	end	else if (num==16'd24623) begin
		isPrime = 1;
	end	else if (num==16'd24631) begin
		isPrime = 1;
	end	else if (num==16'd24659) begin
		isPrime = 1;
	end	else if (num==16'd24671) begin
		isPrime = 1;
	end	else if (num==16'd24677) begin
		isPrime = 1;
	end	else if (num==16'd24683) begin
		isPrime = 1;
	end	else if (num==16'd24691) begin
		isPrime = 1;
	end	else if (num==16'd24697) begin
		isPrime = 1;
	end	else if (num==16'd24709) begin
		isPrime = 1;
	end	else if (num==16'd24733) begin
		isPrime = 1;
	end	else if (num==16'd24749) begin
		isPrime = 1;
	end	else if (num==16'd24763) begin
		isPrime = 1;
	end	else if (num==16'd24767) begin
		isPrime = 1;
	end	else if (num==16'd24781) begin
		isPrime = 1;
	end	else if (num==16'd24793) begin
		isPrime = 1;
	end	else if (num==16'd24799) begin
		isPrime = 1;
	end	else if (num==16'd24809) begin
		isPrime = 1;
	end	else if (num==16'd24821) begin
		isPrime = 1;
	end	else if (num==16'd24841) begin
		isPrime = 1;
	end	else if (num==16'd24847) begin
		isPrime = 1;
	end	else if (num==16'd24851) begin
		isPrime = 1;
	end	else if (num==16'd24859) begin
		isPrime = 1;
	end	else if (num==16'd24877) begin
		isPrime = 1;
	end	else if (num==16'd24889) begin
		isPrime = 1;
	end	else if (num==16'd24907) begin
		isPrime = 1;
	end	else if (num==16'd24917) begin
		isPrime = 1;
	end	else if (num==16'd24919) begin
		isPrime = 1;
	end	else if (num==16'd24923) begin
		isPrime = 1;
	end	else if (num==16'd24943) begin
		isPrime = 1;
	end	else if (num==16'd24953) begin
		isPrime = 1;
	end	else if (num==16'd24967) begin
		isPrime = 1;
	end	else if (num==16'd24971) begin
		isPrime = 1;
	end	else if (num==16'd24977) begin
		isPrime = 1;
	end	else if (num==16'd24979) begin
		isPrime = 1;
	end	else if (num==16'd24989) begin
		isPrime = 1;
	end	else if (num==16'd25013) begin
		isPrime = 1;
	end	else if (num==16'd25031) begin
		isPrime = 1;
	end	else if (num==16'd25033) begin
		isPrime = 1;
	end	else if (num==16'd25037) begin
		isPrime = 1;
	end	else if (num==16'd25057) begin
		isPrime = 1;
	end	else if (num==16'd25073) begin
		isPrime = 1;
	end	else if (num==16'd25087) begin
		isPrime = 1;
	end	else if (num==16'd25097) begin
		isPrime = 1;
	end	else if (num==16'd25111) begin
		isPrime = 1;
	end	else if (num==16'd25117) begin
		isPrime = 1;
	end	else if (num==16'd25121) begin
		isPrime = 1;
	end	else if (num==16'd25127) begin
		isPrime = 1;
	end	else if (num==16'd25147) begin
		isPrime = 1;
	end	else if (num==16'd25153) begin
		isPrime = 1;
	end	else if (num==16'd25163) begin
		isPrime = 1;
	end	else if (num==16'd25169) begin
		isPrime = 1;
	end	else if (num==16'd25171) begin
		isPrime = 1;
	end	else if (num==16'd25183) begin
		isPrime = 1;
	end	else if (num==16'd25189) begin
		isPrime = 1;
	end	else if (num==16'd25219) begin
		isPrime = 1;
	end	else if (num==16'd25229) begin
		isPrime = 1;
	end	else if (num==16'd25237) begin
		isPrime = 1;
	end	else if (num==16'd25243) begin
		isPrime = 1;
	end	else if (num==16'd25247) begin
		isPrime = 1;
	end	else if (num==16'd25253) begin
		isPrime = 1;
	end	else if (num==16'd25261) begin
		isPrime = 1;
	end	else if (num==16'd25301) begin
		isPrime = 1;
	end	else if (num==16'd25303) begin
		isPrime = 1;
	end	else if (num==16'd25307) begin
		isPrime = 1;
	end	else if (num==16'd25309) begin
		isPrime = 1;
	end	else if (num==16'd25321) begin
		isPrime = 1;
	end	else if (num==16'd25339) begin
		isPrime = 1;
	end	else if (num==16'd25343) begin
		isPrime = 1;
	end	else if (num==16'd25349) begin
		isPrime = 1;
	end	else if (num==16'd25357) begin
		isPrime = 1;
	end	else if (num==16'd25367) begin
		isPrime = 1;
	end	else if (num==16'd25373) begin
		isPrime = 1;
	end	else if (num==16'd25391) begin
		isPrime = 1;
	end	else if (num==16'd25409) begin
		isPrime = 1;
	end	else if (num==16'd25411) begin
		isPrime = 1;
	end	else if (num==16'd25423) begin
		isPrime = 1;
	end	else if (num==16'd25439) begin
		isPrime = 1;
	end	else if (num==16'd25447) begin
		isPrime = 1;
	end	else if (num==16'd25453) begin
		isPrime = 1;
	end	else if (num==16'd25457) begin
		isPrime = 1;
	end	else if (num==16'd25463) begin
		isPrime = 1;
	end	else if (num==16'd25469) begin
		isPrime = 1;
	end	else if (num==16'd25471) begin
		isPrime = 1;
	end	else if (num==16'd25523) begin
		isPrime = 1;
	end	else if (num==16'd25537) begin
		isPrime = 1;
	end	else if (num==16'd25541) begin
		isPrime = 1;
	end	else if (num==16'd25561) begin
		isPrime = 1;
	end	else if (num==16'd25577) begin
		isPrime = 1;
	end	else if (num==16'd25579) begin
		isPrime = 1;
	end	else if (num==16'd25583) begin
		isPrime = 1;
	end	else if (num==16'd25589) begin
		isPrime = 1;
	end	else if (num==16'd25601) begin
		isPrime = 1;
	end	else if (num==16'd25603) begin
		isPrime = 1;
	end	else if (num==16'd25609) begin
		isPrime = 1;
	end	else if (num==16'd25621) begin
		isPrime = 1;
	end	else if (num==16'd25633) begin
		isPrime = 1;
	end	else if (num==16'd25639) begin
		isPrime = 1;
	end	else if (num==16'd25643) begin
		isPrime = 1;
	end	else if (num==16'd25657) begin
		isPrime = 1;
	end	else if (num==16'd25667) begin
		isPrime = 1;
	end	else if (num==16'd25673) begin
		isPrime = 1;
	end	else if (num==16'd25679) begin
		isPrime = 1;
	end	else if (num==16'd25693) begin
		isPrime = 1;
	end	else if (num==16'd25703) begin
		isPrime = 1;
	end	else if (num==16'd25717) begin
		isPrime = 1;
	end	else if (num==16'd25733) begin
		isPrime = 1;
	end	else if (num==16'd25741) begin
		isPrime = 1;
	end	else if (num==16'd25747) begin
		isPrime = 1;
	end	else if (num==16'd25759) begin
		isPrime = 1;
	end	else if (num==16'd25763) begin
		isPrime = 1;
	end	else if (num==16'd25771) begin
		isPrime = 1;
	end	else if (num==16'd25793) begin
		isPrime = 1;
	end	else if (num==16'd25799) begin
		isPrime = 1;
	end	else if (num==16'd25801) begin
		isPrime = 1;
	end	else if (num==16'd25819) begin
		isPrime = 1;
	end	else if (num==16'd25841) begin
		isPrime = 1;
	end	else if (num==16'd25847) begin
		isPrime = 1;
	end	else if (num==16'd25849) begin
		isPrime = 1;
	end	else if (num==16'd25867) begin
		isPrime = 1;
	end	else if (num==16'd25873) begin
		isPrime = 1;
	end	else if (num==16'd25889) begin
		isPrime = 1;
	end	else if (num==16'd25903) begin
		isPrime = 1;
	end	else if (num==16'd25913) begin
		isPrime = 1;
	end	else if (num==16'd25919) begin
		isPrime = 1;
	end	else if (num==16'd25931) begin
		isPrime = 1;
	end	else if (num==16'd25933) begin
		isPrime = 1;
	end	else if (num==16'd25939) begin
		isPrime = 1;
	end	else if (num==16'd25943) begin
		isPrime = 1;
	end	else if (num==16'd25951) begin
		isPrime = 1;
	end	else if (num==16'd25969) begin
		isPrime = 1;
	end	else if (num==16'd25981) begin
		isPrime = 1;
	end	else if (num==16'd25997) begin
		isPrime = 1;
	end	else if (num==16'd25999) begin
		isPrime = 1;
	end	else if (num==16'd26003) begin
		isPrime = 1;
	end	else if (num==16'd26017) begin
		isPrime = 1;
	end	else if (num==16'd26021) begin
		isPrime = 1;
	end	else if (num==16'd26029) begin
		isPrime = 1;
	end	else if (num==16'd26041) begin
		isPrime = 1;
	end	else if (num==16'd26053) begin
		isPrime = 1;
	end	else if (num==16'd26083) begin
		isPrime = 1;
	end	else if (num==16'd26099) begin
		isPrime = 1;
	end	else if (num==16'd26107) begin
		isPrime = 1;
	end	else if (num==16'd26111) begin
		isPrime = 1;
	end	else if (num==16'd26113) begin
		isPrime = 1;
	end	else if (num==16'd26119) begin
		isPrime = 1;
	end	else if (num==16'd26141) begin
		isPrime = 1;
	end	else if (num==16'd26153) begin
		isPrime = 1;
	end	else if (num==16'd26161) begin
		isPrime = 1;
	end	else if (num==16'd26171) begin
		isPrime = 1;
	end	else if (num==16'd26177) begin
		isPrime = 1;
	end	else if (num==16'd26183) begin
		isPrime = 1;
	end	else if (num==16'd26189) begin
		isPrime = 1;
	end	else if (num==16'd26203) begin
		isPrime = 1;
	end	else if (num==16'd26209) begin
		isPrime = 1;
	end	else if (num==16'd26227) begin
		isPrime = 1;
	end	else if (num==16'd26237) begin
		isPrime = 1;
	end	else if (num==16'd26249) begin
		isPrime = 1;
	end	else if (num==16'd26251) begin
		isPrime = 1;
	end	else if (num==16'd26261) begin
		isPrime = 1;
	end	else if (num==16'd26263) begin
		isPrime = 1;
	end	else if (num==16'd26267) begin
		isPrime = 1;
	end	else if (num==16'd26293) begin
		isPrime = 1;
	end	else if (num==16'd26297) begin
		isPrime = 1;
	end	else if (num==16'd26309) begin
		isPrime = 1;
	end	else if (num==16'd26317) begin
		isPrime = 1;
	end	else if (num==16'd26321) begin
		isPrime = 1;
	end	else if (num==16'd26339) begin
		isPrime = 1;
	end	else if (num==16'd26347) begin
		isPrime = 1;
	end	else if (num==16'd26357) begin
		isPrime = 1;
	end	else if (num==16'd26371) begin
		isPrime = 1;
	end	else if (num==16'd26387) begin
		isPrime = 1;
	end	else if (num==16'd26393) begin
		isPrime = 1;
	end	else if (num==16'd26399) begin
		isPrime = 1;
	end	else if (num==16'd26407) begin
		isPrime = 1;
	end	else if (num==16'd26417) begin
		isPrime = 1;
	end	else if (num==16'd26423) begin
		isPrime = 1;
	end	else if (num==16'd26431) begin
		isPrime = 1;
	end	else if (num==16'd26437) begin
		isPrime = 1;
	end	else if (num==16'd26449) begin
		isPrime = 1;
	end	else if (num==16'd26459) begin
		isPrime = 1;
	end	else if (num==16'd26479) begin
		isPrime = 1;
	end	else if (num==16'd26489) begin
		isPrime = 1;
	end	else if (num==16'd26497) begin
		isPrime = 1;
	end	else if (num==16'd26501) begin
		isPrime = 1;
	end	else if (num==16'd26513) begin
		isPrime = 1;
	end	else if (num==16'd26539) begin
		isPrime = 1;
	end	else if (num==16'd26557) begin
		isPrime = 1;
	end	else if (num==16'd26561) begin
		isPrime = 1;
	end	else if (num==16'd26573) begin
		isPrime = 1;
	end	else if (num==16'd26591) begin
		isPrime = 1;
	end	else if (num==16'd26597) begin
		isPrime = 1;
	end	else if (num==16'd26627) begin
		isPrime = 1;
	end	else if (num==16'd26633) begin
		isPrime = 1;
	end	else if (num==16'd26641) begin
		isPrime = 1;
	end	else if (num==16'd26647) begin
		isPrime = 1;
	end	else if (num==16'd26669) begin
		isPrime = 1;
	end	else if (num==16'd26681) begin
		isPrime = 1;
	end	else if (num==16'd26683) begin
		isPrime = 1;
	end	else if (num==16'd26687) begin
		isPrime = 1;
	end	else if (num==16'd26693) begin
		isPrime = 1;
	end	else if (num==16'd26699) begin
		isPrime = 1;
	end	else if (num==16'd26701) begin
		isPrime = 1;
	end	else if (num==16'd26711) begin
		isPrime = 1;
	end	else if (num==16'd26713) begin
		isPrime = 1;
	end	else if (num==16'd26717) begin
		isPrime = 1;
	end	else if (num==16'd26723) begin
		isPrime = 1;
	end	else if (num==16'd26729) begin
		isPrime = 1;
	end	else if (num==16'd26731) begin
		isPrime = 1;
	end	else if (num==16'd26737) begin
		isPrime = 1;
	end	else if (num==16'd26759) begin
		isPrime = 1;
	end	else if (num==16'd26777) begin
		isPrime = 1;
	end	else if (num==16'd26783) begin
		isPrime = 1;
	end	else if (num==16'd26801) begin
		isPrime = 1;
	end	else if (num==16'd26813) begin
		isPrime = 1;
	end	else if (num==16'd26821) begin
		isPrime = 1;
	end	else if (num==16'd26833) begin
		isPrime = 1;
	end	else if (num==16'd26839) begin
		isPrime = 1;
	end	else if (num==16'd26849) begin
		isPrime = 1;
	end	else if (num==16'd26861) begin
		isPrime = 1;
	end	else if (num==16'd26863) begin
		isPrime = 1;
	end	else if (num==16'd26879) begin
		isPrime = 1;
	end	else if (num==16'd26881) begin
		isPrime = 1;
	end	else if (num==16'd26891) begin
		isPrime = 1;
	end	else if (num==16'd26893) begin
		isPrime = 1;
	end	else if (num==16'd26903) begin
		isPrime = 1;
	end	else if (num==16'd26921) begin
		isPrime = 1;
	end	else if (num==16'd26927) begin
		isPrime = 1;
	end	else if (num==16'd26947) begin
		isPrime = 1;
	end	else if (num==16'd26951) begin
		isPrime = 1;
	end	else if (num==16'd26953) begin
		isPrime = 1;
	end	else if (num==16'd26959) begin
		isPrime = 1;
	end	else if (num==16'd26981) begin
		isPrime = 1;
	end	else if (num==16'd26987) begin
		isPrime = 1;
	end	else if (num==16'd26993) begin
		isPrime = 1;
	end	else if (num==16'd27011) begin
		isPrime = 1;
	end	else if (num==16'd27017) begin
		isPrime = 1;
	end	else if (num==16'd27031) begin
		isPrime = 1;
	end	else if (num==16'd27043) begin
		isPrime = 1;
	end	else if (num==16'd27059) begin
		isPrime = 1;
	end	else if (num==16'd27061) begin
		isPrime = 1;
	end	else if (num==16'd27067) begin
		isPrime = 1;
	end	else if (num==16'd27073) begin
		isPrime = 1;
	end	else if (num==16'd27077) begin
		isPrime = 1;
	end	else if (num==16'd27091) begin
		isPrime = 1;
	end	else if (num==16'd27103) begin
		isPrime = 1;
	end	else if (num==16'd27107) begin
		isPrime = 1;
	end	else if (num==16'd27109) begin
		isPrime = 1;
	end	else if (num==16'd27127) begin
		isPrime = 1;
	end	else if (num==16'd27143) begin
		isPrime = 1;
	end	else if (num==16'd27179) begin
		isPrime = 1;
	end	else if (num==16'd27191) begin
		isPrime = 1;
	end	else if (num==16'd27197) begin
		isPrime = 1;
	end	else if (num==16'd27211) begin
		isPrime = 1;
	end	else if (num==16'd27239) begin
		isPrime = 1;
	end	else if (num==16'd27241) begin
		isPrime = 1;
	end	else if (num==16'd27253) begin
		isPrime = 1;
	end	else if (num==16'd27259) begin
		isPrime = 1;
	end	else if (num==16'd27271) begin
		isPrime = 1;
	end	else if (num==16'd27277) begin
		isPrime = 1;
	end	else if (num==16'd27281) begin
		isPrime = 1;
	end	else if (num==16'd27283) begin
		isPrime = 1;
	end	else if (num==16'd27299) begin
		isPrime = 1;
	end	else if (num==16'd27329) begin
		isPrime = 1;
	end	else if (num==16'd27337) begin
		isPrime = 1;
	end	else if (num==16'd27361) begin
		isPrime = 1;
	end	else if (num==16'd27367) begin
		isPrime = 1;
	end	else if (num==16'd27397) begin
		isPrime = 1;
	end	else if (num==16'd27407) begin
		isPrime = 1;
	end	else if (num==16'd27409) begin
		isPrime = 1;
	end	else if (num==16'd27427) begin
		isPrime = 1;
	end	else if (num==16'd27431) begin
		isPrime = 1;
	end	else if (num==16'd27437) begin
		isPrime = 1;
	end	else if (num==16'd27449) begin
		isPrime = 1;
	end	else if (num==16'd27457) begin
		isPrime = 1;
	end	else if (num==16'd27479) begin
		isPrime = 1;
	end	else if (num==16'd27481) begin
		isPrime = 1;
	end	else if (num==16'd27487) begin
		isPrime = 1;
	end	else if (num==16'd27509) begin
		isPrime = 1;
	end	else if (num==16'd27527) begin
		isPrime = 1;
	end	else if (num==16'd27529) begin
		isPrime = 1;
	end	else if (num==16'd27539) begin
		isPrime = 1;
	end	else if (num==16'd27541) begin
		isPrime = 1;
	end	else if (num==16'd27551) begin
		isPrime = 1;
	end	else if (num==16'd27581) begin
		isPrime = 1;
	end	else if (num==16'd27583) begin
		isPrime = 1;
	end	else if (num==16'd27611) begin
		isPrime = 1;
	end	else if (num==16'd27617) begin
		isPrime = 1;
	end	else if (num==16'd27631) begin
		isPrime = 1;
	end	else if (num==16'd27647) begin
		isPrime = 1;
	end	else if (num==16'd27653) begin
		isPrime = 1;
	end	else if (num==16'd27673) begin
		isPrime = 1;
	end	else if (num==16'd27689) begin
		isPrime = 1;
	end	else if (num==16'd27691) begin
		isPrime = 1;
	end	else if (num==16'd27697) begin
		isPrime = 1;
	end	else if (num==16'd27701) begin
		isPrime = 1;
	end	else if (num==16'd27733) begin
		isPrime = 1;
	end	else if (num==16'd27737) begin
		isPrime = 1;
	end	else if (num==16'd27739) begin
		isPrime = 1;
	end	else if (num==16'd27743) begin
		isPrime = 1;
	end	else if (num==16'd27749) begin
		isPrime = 1;
	end	else if (num==16'd27751) begin
		isPrime = 1;
	end	else if (num==16'd27763) begin
		isPrime = 1;
	end	else if (num==16'd27767) begin
		isPrime = 1;
	end	else if (num==16'd27773) begin
		isPrime = 1;
	end	else if (num==16'd27779) begin
		isPrime = 1;
	end	else if (num==16'd27791) begin
		isPrime = 1;
	end	else if (num==16'd27793) begin
		isPrime = 1;
	end	else if (num==16'd27799) begin
		isPrime = 1;
	end	else if (num==16'd27803) begin
		isPrime = 1;
	end	else if (num==16'd27809) begin
		isPrime = 1;
	end	else if (num==16'd27817) begin
		isPrime = 1;
	end	else if (num==16'd27823) begin
		isPrime = 1;
	end	else if (num==16'd27827) begin
		isPrime = 1;
	end	else if (num==16'd27847) begin
		isPrime = 1;
	end	else if (num==16'd27851) begin
		isPrime = 1;
	end	else if (num==16'd27883) begin
		isPrime = 1;
	end	else if (num==16'd27893) begin
		isPrime = 1;
	end	else if (num==16'd27901) begin
		isPrime = 1;
	end	else if (num==16'd27917) begin
		isPrime = 1;
	end	else if (num==16'd27919) begin
		isPrime = 1;
	end	else if (num==16'd27941) begin
		isPrime = 1;
	end	else if (num==16'd27943) begin
		isPrime = 1;
	end	else if (num==16'd27947) begin
		isPrime = 1;
	end	else if (num==16'd27953) begin
		isPrime = 1;
	end	else if (num==16'd27961) begin
		isPrime = 1;
	end	else if (num==16'd27967) begin
		isPrime = 1;
	end	else if (num==16'd27983) begin
		isPrime = 1;
	end	else if (num==16'd27997) begin
		isPrime = 1;
	end	else if (num==16'd28001) begin
		isPrime = 1;
	end	else if (num==16'd28019) begin
		isPrime = 1;
	end	else if (num==16'd28027) begin
		isPrime = 1;
	end	else if (num==16'd28031) begin
		isPrime = 1;
	end	else if (num==16'd28051) begin
		isPrime = 1;
	end	else if (num==16'd28057) begin
		isPrime = 1;
	end	else if (num==16'd28069) begin
		isPrime = 1;
	end	else if (num==16'd28081) begin
		isPrime = 1;
	end	else if (num==16'd28087) begin
		isPrime = 1;
	end	else if (num==16'd28097) begin
		isPrime = 1;
	end	else if (num==16'd28099) begin
		isPrime = 1;
	end	else if (num==16'd28109) begin
		isPrime = 1;
	end	else if (num==16'd28111) begin
		isPrime = 1;
	end	else if (num==16'd28123) begin
		isPrime = 1;
	end	else if (num==16'd28151) begin
		isPrime = 1;
	end	else if (num==16'd28163) begin
		isPrime = 1;
	end	else if (num==16'd28181) begin
		isPrime = 1;
	end	else if (num==16'd28183) begin
		isPrime = 1;
	end	else if (num==16'd28201) begin
		isPrime = 1;
	end	else if (num==16'd28211) begin
		isPrime = 1;
	end	else if (num==16'd28219) begin
		isPrime = 1;
	end	else if (num==16'd28229) begin
		isPrime = 1;
	end	else if (num==16'd28277) begin
		isPrime = 1;
	end	else if (num==16'd28279) begin
		isPrime = 1;
	end	else if (num==16'd28283) begin
		isPrime = 1;
	end	else if (num==16'd28289) begin
		isPrime = 1;
	end	else if (num==16'd28297) begin
		isPrime = 1;
	end	else if (num==16'd28307) begin
		isPrime = 1;
	end	else if (num==16'd28309) begin
		isPrime = 1;
	end	else if (num==16'd28319) begin
		isPrime = 1;
	end	else if (num==16'd28349) begin
		isPrime = 1;
	end	else if (num==16'd28351) begin
		isPrime = 1;
	end	else if (num==16'd28387) begin
		isPrime = 1;
	end	else if (num==16'd28393) begin
		isPrime = 1;
	end	else if (num==16'd28403) begin
		isPrime = 1;
	end	else if (num==16'd28409) begin
		isPrime = 1;
	end	else if (num==16'd28411) begin
		isPrime = 1;
	end	else if (num==16'd28429) begin
		isPrime = 1;
	end	else if (num==16'd28433) begin
		isPrime = 1;
	end	else if (num==16'd28439) begin
		isPrime = 1;
	end	else if (num==16'd28447) begin
		isPrime = 1;
	end	else if (num==16'd28463) begin
		isPrime = 1;
	end	else if (num==16'd28477) begin
		isPrime = 1;
	end	else if (num==16'd28493) begin
		isPrime = 1;
	end	else if (num==16'd28499) begin
		isPrime = 1;
	end	else if (num==16'd28513) begin
		isPrime = 1;
	end	else if (num==16'd28517) begin
		isPrime = 1;
	end	else if (num==16'd28537) begin
		isPrime = 1;
	end	else if (num==16'd28541) begin
		isPrime = 1;
	end	else if (num==16'd28547) begin
		isPrime = 1;
	end	else if (num==16'd28549) begin
		isPrime = 1;
	end	else if (num==16'd28559) begin
		isPrime = 1;
	end	else if (num==16'd28571) begin
		isPrime = 1;
	end	else if (num==16'd28573) begin
		isPrime = 1;
	end	else if (num==16'd28579) begin
		isPrime = 1;
	end	else if (num==16'd28591) begin
		isPrime = 1;
	end	else if (num==16'd28597) begin
		isPrime = 1;
	end	else if (num==16'd28603) begin
		isPrime = 1;
	end	else if (num==16'd28607) begin
		isPrime = 1;
	end	else if (num==16'd28619) begin
		isPrime = 1;
	end	else if (num==16'd28621) begin
		isPrime = 1;
	end	else if (num==16'd28627) begin
		isPrime = 1;
	end	else if (num==16'd28631) begin
		isPrime = 1;
	end	else if (num==16'd28643) begin
		isPrime = 1;
	end	else if (num==16'd28649) begin
		isPrime = 1;
	end	else if (num==16'd28657) begin
		isPrime = 1;
	end	else if (num==16'd28661) begin
		isPrime = 1;
	end	else if (num==16'd28663) begin
		isPrime = 1;
	end	else if (num==16'd28669) begin
		isPrime = 1;
	end	else if (num==16'd28687) begin
		isPrime = 1;
	end	else if (num==16'd28697) begin
		isPrime = 1;
	end	else if (num==16'd28703) begin
		isPrime = 1;
	end	else if (num==16'd28711) begin
		isPrime = 1;
	end	else if (num==16'd28723) begin
		isPrime = 1;
	end	else if (num==16'd28729) begin
		isPrime = 1;
	end	else if (num==16'd28751) begin
		isPrime = 1;
	end	else if (num==16'd28753) begin
		isPrime = 1;
	end	else if (num==16'd28759) begin
		isPrime = 1;
	end	else if (num==16'd28771) begin
		isPrime = 1;
	end	else if (num==16'd28789) begin
		isPrime = 1;
	end	else if (num==16'd28793) begin
		isPrime = 1;
	end	else if (num==16'd28807) begin
		isPrime = 1;
	end	else if (num==16'd28813) begin
		isPrime = 1;
	end	else if (num==16'd28817) begin
		isPrime = 1;
	end	else if (num==16'd28837) begin
		isPrime = 1;
	end	else if (num==16'd28843) begin
		isPrime = 1;
	end	else if (num==16'd28859) begin
		isPrime = 1;
	end	else if (num==16'd28867) begin
		isPrime = 1;
	end	else if (num==16'd28871) begin
		isPrime = 1;
	end	else if (num==16'd28879) begin
		isPrime = 1;
	end	else if (num==16'd28901) begin
		isPrime = 1;
	end	else if (num==16'd28909) begin
		isPrime = 1;
	end	else if (num==16'd28921) begin
		isPrime = 1;
	end	else if (num==16'd28927) begin
		isPrime = 1;
	end	else if (num==16'd28933) begin
		isPrime = 1;
	end	else if (num==16'd28949) begin
		isPrime = 1;
	end	else if (num==16'd28961) begin
		isPrime = 1;
	end	else if (num==16'd28979) begin
		isPrime = 1;
	end	else if (num==16'd29009) begin
		isPrime = 1;
	end	else if (num==16'd29017) begin
		isPrime = 1;
	end	else if (num==16'd29021) begin
		isPrime = 1;
	end	else if (num==16'd29023) begin
		isPrime = 1;
	end	else if (num==16'd29027) begin
		isPrime = 1;
	end	else if (num==16'd29033) begin
		isPrime = 1;
	end	else if (num==16'd29059) begin
		isPrime = 1;
	end	else if (num==16'd29063) begin
		isPrime = 1;
	end	else if (num==16'd29077) begin
		isPrime = 1;
	end	else if (num==16'd29101) begin
		isPrime = 1;
	end	else if (num==16'd29123) begin
		isPrime = 1;
	end	else if (num==16'd29129) begin
		isPrime = 1;
	end	else if (num==16'd29131) begin
		isPrime = 1;
	end	else if (num==16'd29137) begin
		isPrime = 1;
	end	else if (num==16'd29147) begin
		isPrime = 1;
	end	else if (num==16'd29153) begin
		isPrime = 1;
	end	else if (num==16'd29167) begin
		isPrime = 1;
	end	else if (num==16'd29173) begin
		isPrime = 1;
	end	else if (num==16'd29179) begin
		isPrime = 1;
	end	else if (num==16'd29191) begin
		isPrime = 1;
	end	else if (num==16'd29201) begin
		isPrime = 1;
	end	else if (num==16'd29207) begin
		isPrime = 1;
	end	else if (num==16'd29209) begin
		isPrime = 1;
	end	else if (num==16'd29221) begin
		isPrime = 1;
	end	else if (num==16'd29231) begin
		isPrime = 1;
	end	else if (num==16'd29243) begin
		isPrime = 1;
	end	else if (num==16'd29251) begin
		isPrime = 1;
	end	else if (num==16'd29269) begin
		isPrime = 1;
	end	else if (num==16'd29287) begin
		isPrime = 1;
	end	else if (num==16'd29297) begin
		isPrime = 1;
	end	else if (num==16'd29303) begin
		isPrime = 1;
	end	else if (num==16'd29311) begin
		isPrime = 1;
	end	else if (num==16'd29327) begin
		isPrime = 1;
	end	else if (num==16'd29333) begin
		isPrime = 1;
	end	else if (num==16'd29339) begin
		isPrime = 1;
	end	else if (num==16'd29347) begin
		isPrime = 1;
	end	else if (num==16'd29363) begin
		isPrime = 1;
	end	else if (num==16'd29383) begin
		isPrime = 1;
	end	else if (num==16'd29387) begin
		isPrime = 1;
	end	else if (num==16'd29389) begin
		isPrime = 1;
	end	else if (num==16'd29399) begin
		isPrime = 1;
	end	else if (num==16'd29401) begin
		isPrime = 1;
	end	else if (num==16'd29411) begin
		isPrime = 1;
	end	else if (num==16'd29423) begin
		isPrime = 1;
	end	else if (num==16'd29429) begin
		isPrime = 1;
	end	else if (num==16'd29437) begin
		isPrime = 1;
	end	else if (num==16'd29443) begin
		isPrime = 1;
	end	else if (num==16'd29453) begin
		isPrime = 1;
	end	else if (num==16'd29473) begin
		isPrime = 1;
	end	else if (num==16'd29483) begin
		isPrime = 1;
	end	else if (num==16'd29501) begin
		isPrime = 1;
	end	else if (num==16'd29527) begin
		isPrime = 1;
	end	else if (num==16'd29531) begin
		isPrime = 1;
	end	else if (num==16'd29537) begin
		isPrime = 1;
	end	else if (num==16'd29567) begin
		isPrime = 1;
	end	else if (num==16'd29569) begin
		isPrime = 1;
	end	else if (num==16'd29573) begin
		isPrime = 1;
	end	else if (num==16'd29581) begin
		isPrime = 1;
	end	else if (num==16'd29587) begin
		isPrime = 1;
	end	else if (num==16'd29599) begin
		isPrime = 1;
	end	else if (num==16'd29611) begin
		isPrime = 1;
	end	else if (num==16'd29629) begin
		isPrime = 1;
	end	else if (num==16'd29633) begin
		isPrime = 1;
	end	else if (num==16'd29641) begin
		isPrime = 1;
	end	else if (num==16'd29663) begin
		isPrime = 1;
	end	else if (num==16'd29669) begin
		isPrime = 1;
	end	else if (num==16'd29671) begin
		isPrime = 1;
	end	else if (num==16'd29683) begin
		isPrime = 1;
	end	else if (num==16'd29717) begin
		isPrime = 1;
	end	else if (num==16'd29723) begin
		isPrime = 1;
	end	else if (num==16'd29741) begin
		isPrime = 1;
	end	else if (num==16'd29753) begin
		isPrime = 1;
	end	else if (num==16'd29759) begin
		isPrime = 1;
	end	else if (num==16'd29761) begin
		isPrime = 1;
	end	else if (num==16'd29789) begin
		isPrime = 1;
	end	else if (num==16'd29803) begin
		isPrime = 1;
	end	else if (num==16'd29819) begin
		isPrime = 1;
	end	else if (num==16'd29833) begin
		isPrime = 1;
	end	else if (num==16'd29837) begin
		isPrime = 1;
	end	else if (num==16'd29851) begin
		isPrime = 1;
	end	else if (num==16'd29863) begin
		isPrime = 1;
	end	else if (num==16'd29867) begin
		isPrime = 1;
	end	else if (num==16'd29873) begin
		isPrime = 1;
	end	else if (num==16'd29879) begin
		isPrime = 1;
	end	else if (num==16'd29881) begin
		isPrime = 1;
	end	else if (num==16'd29917) begin
		isPrime = 1;
	end	else if (num==16'd29921) begin
		isPrime = 1;
	end	else if (num==16'd29927) begin
		isPrime = 1;
	end	else if (num==16'd29947) begin
		isPrime = 1;
	end	else if (num==16'd29959) begin
		isPrime = 1;
	end	else if (num==16'd29983) begin
		isPrime = 1;
	end	else if (num==16'd29989) begin
		isPrime = 1;
	end	else if (num==16'd30011) begin
		isPrime = 1;
	end	else if (num==16'd30013) begin
		isPrime = 1;
	end	else if (num==16'd30029) begin
		isPrime = 1;
	end	else if (num==16'd30047) begin
		isPrime = 1;
	end	else if (num==16'd30059) begin
		isPrime = 1;
	end	else if (num==16'd30071) begin
		isPrime = 1;
	end	else if (num==16'd30089) begin
		isPrime = 1;
	end	else if (num==16'd30091) begin
		isPrime = 1;
	end	else if (num==16'd30097) begin
		isPrime = 1;
	end	else if (num==16'd30103) begin
		isPrime = 1;
	end	else if (num==16'd30109) begin
		isPrime = 1;
	end	else if (num==16'd30113) begin
		isPrime = 1;
	end	else if (num==16'd30119) begin
		isPrime = 1;
	end	else if (num==16'd30133) begin
		isPrime = 1;
	end	else if (num==16'd30137) begin
		isPrime = 1;
	end	else if (num==16'd30139) begin
		isPrime = 1;
	end	else if (num==16'd30161) begin
		isPrime = 1;
	end	else if (num==16'd30169) begin
		isPrime = 1;
	end	else if (num==16'd30181) begin
		isPrime = 1;
	end	else if (num==16'd30187) begin
		isPrime = 1;
	end	else if (num==16'd30197) begin
		isPrime = 1;
	end	else if (num==16'd30203) begin
		isPrime = 1;
	end	else if (num==16'd30211) begin
		isPrime = 1;
	end	else if (num==16'd30223) begin
		isPrime = 1;
	end	else if (num==16'd30241) begin
		isPrime = 1;
	end	else if (num==16'd30253) begin
		isPrime = 1;
	end	else if (num==16'd30259) begin
		isPrime = 1;
	end	else if (num==16'd30269) begin
		isPrime = 1;
	end	else if (num==16'd30271) begin
		isPrime = 1;
	end	else if (num==16'd30293) begin
		isPrime = 1;
	end	else if (num==16'd30307) begin
		isPrime = 1;
	end	else if (num==16'd30313) begin
		isPrime = 1;
	end	else if (num==16'd30319) begin
		isPrime = 1;
	end	else if (num==16'd30323) begin
		isPrime = 1;
	end	else if (num==16'd30341) begin
		isPrime = 1;
	end	else if (num==16'd30347) begin
		isPrime = 1;
	end	else if (num==16'd30367) begin
		isPrime = 1;
	end	else if (num==16'd30389) begin
		isPrime = 1;
	end	else if (num==16'd30391) begin
		isPrime = 1;
	end	else if (num==16'd30403) begin
		isPrime = 1;
	end	else if (num==16'd30427) begin
		isPrime = 1;
	end	else if (num==16'd30431) begin
		isPrime = 1;
	end	else if (num==16'd30449) begin
		isPrime = 1;
	end	else if (num==16'd30467) begin
		isPrime = 1;
	end	else if (num==16'd30469) begin
		isPrime = 1;
	end	else if (num==16'd30491) begin
		isPrime = 1;
	end	else if (num==16'd30493) begin
		isPrime = 1;
	end	else if (num==16'd30497) begin
		isPrime = 1;
	end	else if (num==16'd30509) begin
		isPrime = 1;
	end	else if (num==16'd30517) begin
		isPrime = 1;
	end	else if (num==16'd30529) begin
		isPrime = 1;
	end	else if (num==16'd30539) begin
		isPrime = 1;
	end	else if (num==16'd30553) begin
		isPrime = 1;
	end	else if (num==16'd30557) begin
		isPrime = 1;
	end	else if (num==16'd30559) begin
		isPrime = 1;
	end	else if (num==16'd30577) begin
		isPrime = 1;
	end	else if (num==16'd30593) begin
		isPrime = 1;
	end	else if (num==16'd30631) begin
		isPrime = 1;
	end	else if (num==16'd30637) begin
		isPrime = 1;
	end	else if (num==16'd30643) begin
		isPrime = 1;
	end	else if (num==16'd30649) begin
		isPrime = 1;
	end	else if (num==16'd30661) begin
		isPrime = 1;
	end	else if (num==16'd30671) begin
		isPrime = 1;
	end	else if (num==16'd30677) begin
		isPrime = 1;
	end	else if (num==16'd30689) begin
		isPrime = 1;
	end	else if (num==16'd30697) begin
		isPrime = 1;
	end	else if (num==16'd30703) begin
		isPrime = 1;
	end	else if (num==16'd30707) begin
		isPrime = 1;
	end	else if (num==16'd30713) begin
		isPrime = 1;
	end	else if (num==16'd30727) begin
		isPrime = 1;
	end	else if (num==16'd30757) begin
		isPrime = 1;
	end	else if (num==16'd30763) begin
		isPrime = 1;
	end	else if (num==16'd30773) begin
		isPrime = 1;
	end	else if (num==16'd30781) begin
		isPrime = 1;
	end	else if (num==16'd30803) begin
		isPrime = 1;
	end	else if (num==16'd30809) begin
		isPrime = 1;
	end	else if (num==16'd30817) begin
		isPrime = 1;
	end	else if (num==16'd30829) begin
		isPrime = 1;
	end	else if (num==16'd30839) begin
		isPrime = 1;
	end	else if (num==16'd30841) begin
		isPrime = 1;
	end	else if (num==16'd30851) begin
		isPrime = 1;
	end	else if (num==16'd30853) begin
		isPrime = 1;
	end	else if (num==16'd30859) begin
		isPrime = 1;
	end	else if (num==16'd30869) begin
		isPrime = 1;
	end	else if (num==16'd30871) begin
		isPrime = 1;
	end	else if (num==16'd30881) begin
		isPrime = 1;
	end	else if (num==16'd30893) begin
		isPrime = 1;
	end	else if (num==16'd30911) begin
		isPrime = 1;
	end	else if (num==16'd30931) begin
		isPrime = 1;
	end	else if (num==16'd30937) begin
		isPrime = 1;
	end	else if (num==16'd30941) begin
		isPrime = 1;
	end	else if (num==16'd30949) begin
		isPrime = 1;
	end	else if (num==16'd30971) begin
		isPrime = 1;
	end	else if (num==16'd30977) begin
		isPrime = 1;
	end	else if (num==16'd30983) begin
		isPrime = 1;
	end	else if (num==16'd31013) begin
		isPrime = 1;
	end	else if (num==16'd31019) begin
		isPrime = 1;
	end	else if (num==16'd31033) begin
		isPrime = 1;
	end	else if (num==16'd31039) begin
		isPrime = 1;
	end	else if (num==16'd31051) begin
		isPrime = 1;
	end	else if (num==16'd31063) begin
		isPrime = 1;
	end	else if (num==16'd31069) begin
		isPrime = 1;
	end	else if (num==16'd31079) begin
		isPrime = 1;
	end	else if (num==16'd31081) begin
		isPrime = 1;
	end	else if (num==16'd31091) begin
		isPrime = 1;
	end	else if (num==16'd31121) begin
		isPrime = 1;
	end	else if (num==16'd31123) begin
		isPrime = 1;
	end	else if (num==16'd31139) begin
		isPrime = 1;
	end	else if (num==16'd31147) begin
		isPrime = 1;
	end	else if (num==16'd31151) begin
		isPrime = 1;
	end	else if (num==16'd31153) begin
		isPrime = 1;
	end	else if (num==16'd31159) begin
		isPrime = 1;
	end	else if (num==16'd31177) begin
		isPrime = 1;
	end	else if (num==16'd31181) begin
		isPrime = 1;
	end	else if (num==16'd31183) begin
		isPrime = 1;
	end	else if (num==16'd31189) begin
		isPrime = 1;
	end	else if (num==16'd31193) begin
		isPrime = 1;
	end	else if (num==16'd31219) begin
		isPrime = 1;
	end	else if (num==16'd31223) begin
		isPrime = 1;
	end	else if (num==16'd31231) begin
		isPrime = 1;
	end	else if (num==16'd31237) begin
		isPrime = 1;
	end	else if (num==16'd31247) begin
		isPrime = 1;
	end	else if (num==16'd31249) begin
		isPrime = 1;
	end	else if (num==16'd31253) begin
		isPrime = 1;
	end	else if (num==16'd31259) begin
		isPrime = 1;
	end	else if (num==16'd31267) begin
		isPrime = 1;
	end	else if (num==16'd31271) begin
		isPrime = 1;
	end	else if (num==16'd31277) begin
		isPrime = 1;
	end	else if (num==16'd31307) begin
		isPrime = 1;
	end	else if (num==16'd31319) begin
		isPrime = 1;
	end	else if (num==16'd31321) begin
		isPrime = 1;
	end	else if (num==16'd31327) begin
		isPrime = 1;
	end	else if (num==16'd31333) begin
		isPrime = 1;
	end	else if (num==16'd31337) begin
		isPrime = 1;
	end	else if (num==16'd31357) begin
		isPrime = 1;
	end	else if (num==16'd31379) begin
		isPrime = 1;
	end	else if (num==16'd31387) begin
		isPrime = 1;
	end	else if (num==16'd31391) begin
		isPrime = 1;
	end	else if (num==16'd31393) begin
		isPrime = 1;
	end	else if (num==16'd31397) begin
		isPrime = 1;
	end	else if (num==16'd31469) begin
		isPrime = 1;
	end	else if (num==16'd31477) begin
		isPrime = 1;
	end	else if (num==16'd31481) begin
		isPrime = 1;
	end	else if (num==16'd31489) begin
		isPrime = 1;
	end	else if (num==16'd31511) begin
		isPrime = 1;
	end	else if (num==16'd31513) begin
		isPrime = 1;
	end	else if (num==16'd31517) begin
		isPrime = 1;
	end	else if (num==16'd31531) begin
		isPrime = 1;
	end	else if (num==16'd31541) begin
		isPrime = 1;
	end	else if (num==16'd31543) begin
		isPrime = 1;
	end	else if (num==16'd31547) begin
		isPrime = 1;
	end	else if (num==16'd31567) begin
		isPrime = 1;
	end	else if (num==16'd31573) begin
		isPrime = 1;
	end	else if (num==16'd31583) begin
		isPrime = 1;
	end	else if (num==16'd31601) begin
		isPrime = 1;
	end	else if (num==16'd31607) begin
		isPrime = 1;
	end	else if (num==16'd31627) begin
		isPrime = 1;
	end	else if (num==16'd31643) begin
		isPrime = 1;
	end	else if (num==16'd31649) begin
		isPrime = 1;
	end	else if (num==16'd31657) begin
		isPrime = 1;
	end	else if (num==16'd31663) begin
		isPrime = 1;
	end	else if (num==16'd31667) begin
		isPrime = 1;
	end	else if (num==16'd31687) begin
		isPrime = 1;
	end	else if (num==16'd31699) begin
		isPrime = 1;
	end	else if (num==16'd31721) begin
		isPrime = 1;
	end	else if (num==16'd31723) begin
		isPrime = 1;
	end	else if (num==16'd31727) begin
		isPrime = 1;
	end	else if (num==16'd31729) begin
		isPrime = 1;
	end	else if (num==16'd31741) begin
		isPrime = 1;
	end	else if (num==16'd31751) begin
		isPrime = 1;
	end	else if (num==16'd31769) begin
		isPrime = 1;
	end	else if (num==16'd31771) begin
		isPrime = 1;
	end	else if (num==16'd31793) begin
		isPrime = 1;
	end	else if (num==16'd31799) begin
		isPrime = 1;
	end	else if (num==16'd31817) begin
		isPrime = 1;
	end	else if (num==16'd31847) begin
		isPrime = 1;
	end	else if (num==16'd31849) begin
		isPrime = 1;
	end	else if (num==16'd31859) begin
		isPrime = 1;
	end	else if (num==16'd31873) begin
		isPrime = 1;
	end	else if (num==16'd31883) begin
		isPrime = 1;
	end	else if (num==16'd31891) begin
		isPrime = 1;
	end	else if (num==16'd31907) begin
		isPrime = 1;
	end	else if (num==16'd31957) begin
		isPrime = 1;
	end	else if (num==16'd31963) begin
		isPrime = 1;
	end	else if (num==16'd31973) begin
		isPrime = 1;
	end	else if (num==16'd31981) begin
		isPrime = 1;
	end	else if (num==16'd31991) begin
		isPrime = 1;
	end	else if (num==16'd32003) begin
		isPrime = 1;
	end	else if (num==16'd32009) begin
		isPrime = 1;
	end	else if (num==16'd32027) begin
		isPrime = 1;
	end	else if (num==16'd32029) begin
		isPrime = 1;
	end	else if (num==16'd32051) begin
		isPrime = 1;
	end	else if (num==16'd32057) begin
		isPrime = 1;
	end	else if (num==16'd32059) begin
		isPrime = 1;
	end	else if (num==16'd32063) begin
		isPrime = 1;
	end	else if (num==16'd32069) begin
		isPrime = 1;
	end	else if (num==16'd32077) begin
		isPrime = 1;
	end	else if (num==16'd32083) begin
		isPrime = 1;
	end	else if (num==16'd32089) begin
		isPrime = 1;
	end	else if (num==16'd32099) begin
		isPrime = 1;
	end	else if (num==16'd32117) begin
		isPrime = 1;
	end	else if (num==16'd32119) begin
		isPrime = 1;
	end	else if (num==16'd32141) begin
		isPrime = 1;
	end	else if (num==16'd32143) begin
		isPrime = 1;
	end	else if (num==16'd32159) begin
		isPrime = 1;
	end	else if (num==16'd32173) begin
		isPrime = 1;
	end	else if (num==16'd32183) begin
		isPrime = 1;
	end	else if (num==16'd32189) begin
		isPrime = 1;
	end	else if (num==16'd32191) begin
		isPrime = 1;
	end	else if (num==16'd32203) begin
		isPrime = 1;
	end	else if (num==16'd32213) begin
		isPrime = 1;
	end	else if (num==16'd32233) begin
		isPrime = 1;
	end	else if (num==16'd32237) begin
		isPrime = 1;
	end	else if (num==16'd32251) begin
		isPrime = 1;
	end	else if (num==16'd32257) begin
		isPrime = 1;
	end	else if (num==16'd32261) begin
		isPrime = 1;
	end	else if (num==16'd32297) begin
		isPrime = 1;
	end	else if (num==16'd32299) begin
		isPrime = 1;
	end	else if (num==16'd32303) begin
		isPrime = 1;
	end	else if (num==16'd32309) begin
		isPrime = 1;
	end	else if (num==16'd32321) begin
		isPrime = 1;
	end	else if (num==16'd32323) begin
		isPrime = 1;
	end	else if (num==16'd32327) begin
		isPrime = 1;
	end	else if (num==16'd32341) begin
		isPrime = 1;
	end	else if (num==16'd32353) begin
		isPrime = 1;
	end	else if (num==16'd32359) begin
		isPrime = 1;
	end	else if (num==16'd32363) begin
		isPrime = 1;
	end	else if (num==16'd32369) begin
		isPrime = 1;
	end	else if (num==16'd32371) begin
		isPrime = 1;
	end	else if (num==16'd32377) begin
		isPrime = 1;
	end	else if (num==16'd32381) begin
		isPrime = 1;
	end	else if (num==16'd32401) begin
		isPrime = 1;
	end	else if (num==16'd32411) begin
		isPrime = 1;
	end	else if (num==16'd32413) begin
		isPrime = 1;
	end	else if (num==16'd32423) begin
		isPrime = 1;
	end	else if (num==16'd32429) begin
		isPrime = 1;
	end	else if (num==16'd32441) begin
		isPrime = 1;
	end	else if (num==16'd32443) begin
		isPrime = 1;
	end	else if (num==16'd32467) begin
		isPrime = 1;
	end	else if (num==16'd32479) begin
		isPrime = 1;
	end	else if (num==16'd32491) begin
		isPrime = 1;
	end	else if (num==16'd32497) begin
		isPrime = 1;
	end	else if (num==16'd32503) begin
		isPrime = 1;
	end	else if (num==16'd32507) begin
		isPrime = 1;
	end	else if (num==16'd32531) begin
		isPrime = 1;
	end	else if (num==16'd32533) begin
		isPrime = 1;
	end	else if (num==16'd32537) begin
		isPrime = 1;
	end	else if (num==16'd32561) begin
		isPrime = 1;
	end	else if (num==16'd32563) begin
		isPrime = 1;
	end	else if (num==16'd32569) begin
		isPrime = 1;
	end	else if (num==16'd32573) begin
		isPrime = 1;
	end	else if (num==16'd32579) begin
		isPrime = 1;
	end	else if (num==16'd32587) begin
		isPrime = 1;
	end	else if (num==16'd32603) begin
		isPrime = 1;
	end	else if (num==16'd32609) begin
		isPrime = 1;
	end	else if (num==16'd32611) begin
		isPrime = 1;
	end	else if (num==16'd32621) begin
		isPrime = 1;
	end	else if (num==16'd32633) begin
		isPrime = 1;
	end	else if (num==16'd32647) begin
		isPrime = 1;
	end	else if (num==16'd32653) begin
		isPrime = 1;
	end	else if (num==16'd32687) begin
		isPrime = 1;
	end	else if (num==16'd32693) begin
		isPrime = 1;
	end	else if (num==16'd32707) begin
		isPrime = 1;
	end	else if (num==16'd32713) begin
		isPrime = 1;
	end	else if (num==16'd32717) begin
		isPrime = 1;
	end	else if (num==16'd32719) begin
		isPrime = 1;
	end	else if (num==16'd32749) begin
		isPrime = 1;
	end	else if (num==16'd32771) begin
		isPrime = 1;
	end	else if (num==16'd32779) begin
		isPrime = 1;
	end	else if (num==16'd32783) begin
		isPrime = 1;
	end	else if (num==16'd32789) begin
		isPrime = 1;
	end	else if (num==16'd32797) begin
		isPrime = 1;
	end	else if (num==16'd32801) begin
		isPrime = 1;
	end	else if (num==16'd32803) begin
		isPrime = 1;
	end	else if (num==16'd32831) begin
		isPrime = 1;
	end	else if (num==16'd32833) begin
		isPrime = 1;
	end	else if (num==16'd32839) begin
		isPrime = 1;
	end	else if (num==16'd32843) begin
		isPrime = 1;
	end	else if (num==16'd32869) begin
		isPrime = 1;
	end	else if (num==16'd32887) begin
		isPrime = 1;
	end	else if (num==16'd32909) begin
		isPrime = 1;
	end	else if (num==16'd32911) begin
		isPrime = 1;
	end	else if (num==16'd32917) begin
		isPrime = 1;
	end	else if (num==16'd32933) begin
		isPrime = 1;
	end	else if (num==16'd32939) begin
		isPrime = 1;
	end	else if (num==16'd32941) begin
		isPrime = 1;
	end	else if (num==16'd32957) begin
		isPrime = 1;
	end	else if (num==16'd32969) begin
		isPrime = 1;
	end	else if (num==16'd32971) begin
		isPrime = 1;
	end	else if (num==16'd32983) begin
		isPrime = 1;
	end	else if (num==16'd32987) begin
		isPrime = 1;
	end	else if (num==16'd32993) begin
		isPrime = 1;
	end	else if (num==16'd32999) begin
		isPrime = 1;
	end	else if (num==16'd33013) begin
		isPrime = 1;
	end	else if (num==16'd33023) begin
		isPrime = 1;
	end	else if (num==16'd33029) begin
		isPrime = 1;
	end	else if (num==16'd33037) begin
		isPrime = 1;
	end	else if (num==16'd33049) begin
		isPrime = 1;
	end	else if (num==16'd33053) begin
		isPrime = 1;
	end	else if (num==16'd33071) begin
		isPrime = 1;
	end	else if (num==16'd33073) begin
		isPrime = 1;
	end	else if (num==16'd33083) begin
		isPrime = 1;
	end	else if (num==16'd33091) begin
		isPrime = 1;
	end	else if (num==16'd33107) begin
		isPrime = 1;
	end	else if (num==16'd33113) begin
		isPrime = 1;
	end	else if (num==16'd33119) begin
		isPrime = 1;
	end	else if (num==16'd33149) begin
		isPrime = 1;
	end	else if (num==16'd33151) begin
		isPrime = 1;
	end	else if (num==16'd33161) begin
		isPrime = 1;
	end	else if (num==16'd33179) begin
		isPrime = 1;
	end	else if (num==16'd33181) begin
		isPrime = 1;
	end	else if (num==16'd33191) begin
		isPrime = 1;
	end	else if (num==16'd33199) begin
		isPrime = 1;
	end	else if (num==16'd33203) begin
		isPrime = 1;
	end	else if (num==16'd33211) begin
		isPrime = 1;
	end	else if (num==16'd33223) begin
		isPrime = 1;
	end	else if (num==16'd33247) begin
		isPrime = 1;
	end	else if (num==16'd33287) begin
		isPrime = 1;
	end	else if (num==16'd33289) begin
		isPrime = 1;
	end	else if (num==16'd33301) begin
		isPrime = 1;
	end	else if (num==16'd33311) begin
		isPrime = 1;
	end	else if (num==16'd33317) begin
		isPrime = 1;
	end	else if (num==16'd33329) begin
		isPrime = 1;
	end	else if (num==16'd33331) begin
		isPrime = 1;
	end	else if (num==16'd33343) begin
		isPrime = 1;
	end	else if (num==16'd33347) begin
		isPrime = 1;
	end	else if (num==16'd33349) begin
		isPrime = 1;
	end	else if (num==16'd33353) begin
		isPrime = 1;
	end	else if (num==16'd33359) begin
		isPrime = 1;
	end	else if (num==16'd33377) begin
		isPrime = 1;
	end	else if (num==16'd33391) begin
		isPrime = 1;
	end	else if (num==16'd33403) begin
		isPrime = 1;
	end	else if (num==16'd33409) begin
		isPrime = 1;
	end	else if (num==16'd33413) begin
		isPrime = 1;
	end	else if (num==16'd33427) begin
		isPrime = 1;
	end	else if (num==16'd33457) begin
		isPrime = 1;
	end	else if (num==16'd33461) begin
		isPrime = 1;
	end	else if (num==16'd33469) begin
		isPrime = 1;
	end	else if (num==16'd33479) begin
		isPrime = 1;
	end	else if (num==16'd33487) begin
		isPrime = 1;
	end	else if (num==16'd33493) begin
		isPrime = 1;
	end	else if (num==16'd33503) begin
		isPrime = 1;
	end	else if (num==16'd33521) begin
		isPrime = 1;
	end	else if (num==16'd33529) begin
		isPrime = 1;
	end	else if (num==16'd33533) begin
		isPrime = 1;
	end	else if (num==16'd33547) begin
		isPrime = 1;
	end	else if (num==16'd33563) begin
		isPrime = 1;
	end	else if (num==16'd33569) begin
		isPrime = 1;
	end	else if (num==16'd33577) begin
		isPrime = 1;
	end	else if (num==16'd33581) begin
		isPrime = 1;
	end	else if (num==16'd33587) begin
		isPrime = 1;
	end	else if (num==16'd33589) begin
		isPrime = 1;
	end	else if (num==16'd33599) begin
		isPrime = 1;
	end	else if (num==16'd33601) begin
		isPrime = 1;
	end	else if (num==16'd33613) begin
		isPrime = 1;
	end	else if (num==16'd33617) begin
		isPrime = 1;
	end	else if (num==16'd33619) begin
		isPrime = 1;
	end	else if (num==16'd33623) begin
		isPrime = 1;
	end	else if (num==16'd33629) begin
		isPrime = 1;
	end	else if (num==16'd33637) begin
		isPrime = 1;
	end	else if (num==16'd33641) begin
		isPrime = 1;
	end	else if (num==16'd33647) begin
		isPrime = 1;
	end	else if (num==16'd33679) begin
		isPrime = 1;
	end	else if (num==16'd33703) begin
		isPrime = 1;
	end	else if (num==16'd33713) begin
		isPrime = 1;
	end	else if (num==16'd33721) begin
		isPrime = 1;
	end	else if (num==16'd33739) begin
		isPrime = 1;
	end	else if (num==16'd33749) begin
		isPrime = 1;
	end	else if (num==16'd33751) begin
		isPrime = 1;
	end	else if (num==16'd33757) begin
		isPrime = 1;
	end	else if (num==16'd33767) begin
		isPrime = 1;
	end	else if (num==16'd33769) begin
		isPrime = 1;
	end	else if (num==16'd33773) begin
		isPrime = 1;
	end	else if (num==16'd33791) begin
		isPrime = 1;
	end	else if (num==16'd33797) begin
		isPrime = 1;
	end	else if (num==16'd33809) begin
		isPrime = 1;
	end	else if (num==16'd33811) begin
		isPrime = 1;
	end	else if (num==16'd33827) begin
		isPrime = 1;
	end	else if (num==16'd33829) begin
		isPrime = 1;
	end	else if (num==16'd33851) begin
		isPrime = 1;
	end	else if (num==16'd33857) begin
		isPrime = 1;
	end	else if (num==16'd33863) begin
		isPrime = 1;
	end	else if (num==16'd33871) begin
		isPrime = 1;
	end	else if (num==16'd33889) begin
		isPrime = 1;
	end	else if (num==16'd33893) begin
		isPrime = 1;
	end	else if (num==16'd33911) begin
		isPrime = 1;
	end	else if (num==16'd33923) begin
		isPrime = 1;
	end	else if (num==16'd33931) begin
		isPrime = 1;
	end	else if (num==16'd33937) begin
		isPrime = 1;
	end	else if (num==16'd33941) begin
		isPrime = 1;
	end	else if (num==16'd33961) begin
		isPrime = 1;
	end	else if (num==16'd33967) begin
		isPrime = 1;
	end	else if (num==16'd33997) begin
		isPrime = 1;
	end	else if (num==16'd34019) begin
		isPrime = 1;
	end	else if (num==16'd34031) begin
		isPrime = 1;
	end	else if (num==16'd34033) begin
		isPrime = 1;
	end	else if (num==16'd34039) begin
		isPrime = 1;
	end	else if (num==16'd34057) begin
		isPrime = 1;
	end	else if (num==16'd34061) begin
		isPrime = 1;
	end	else if (num==16'd34123) begin
		isPrime = 1;
	end	else if (num==16'd34127) begin
		isPrime = 1;
	end	else if (num==16'd34129) begin
		isPrime = 1;
	end	else if (num==16'd34141) begin
		isPrime = 1;
	end	else if (num==16'd34147) begin
		isPrime = 1;
	end	else if (num==16'd34157) begin
		isPrime = 1;
	end	else if (num==16'd34159) begin
		isPrime = 1;
	end	else if (num==16'd34171) begin
		isPrime = 1;
	end	else if (num==16'd34183) begin
		isPrime = 1;
	end	else if (num==16'd34211) begin
		isPrime = 1;
	end	else if (num==16'd34213) begin
		isPrime = 1;
	end	else if (num==16'd34217) begin
		isPrime = 1;
	end	else if (num==16'd34231) begin
		isPrime = 1;
	end	else if (num==16'd34253) begin
		isPrime = 1;
	end	else if (num==16'd34259) begin
		isPrime = 1;
	end	else if (num==16'd34261) begin
		isPrime = 1;
	end	else if (num==16'd34267) begin
		isPrime = 1;
	end	else if (num==16'd34273) begin
		isPrime = 1;
	end	else if (num==16'd34283) begin
		isPrime = 1;
	end	else if (num==16'd34297) begin
		isPrime = 1;
	end	else if (num==16'd34301) begin
		isPrime = 1;
	end	else if (num==16'd34303) begin
		isPrime = 1;
	end	else if (num==16'd34313) begin
		isPrime = 1;
	end	else if (num==16'd34319) begin
		isPrime = 1;
	end	else if (num==16'd34327) begin
		isPrime = 1;
	end	else if (num==16'd34337) begin
		isPrime = 1;
	end	else if (num==16'd34351) begin
		isPrime = 1;
	end	else if (num==16'd34361) begin
		isPrime = 1;
	end	else if (num==16'd34367) begin
		isPrime = 1;
	end	else if (num==16'd34369) begin
		isPrime = 1;
	end	else if (num==16'd34381) begin
		isPrime = 1;
	end	else if (num==16'd34403) begin
		isPrime = 1;
	end	else if (num==16'd34421) begin
		isPrime = 1;
	end	else if (num==16'd34429) begin
		isPrime = 1;
	end	else if (num==16'd34439) begin
		isPrime = 1;
	end	else if (num==16'd34457) begin
		isPrime = 1;
	end	else if (num==16'd34469) begin
		isPrime = 1;
	end	else if (num==16'd34471) begin
		isPrime = 1;
	end	else if (num==16'd34483) begin
		isPrime = 1;
	end	else if (num==16'd34487) begin
		isPrime = 1;
	end	else if (num==16'd34499) begin
		isPrime = 1;
	end	else if (num==16'd34501) begin
		isPrime = 1;
	end	else if (num==16'd34511) begin
		isPrime = 1;
	end	else if (num==16'd34513) begin
		isPrime = 1;
	end	else if (num==16'd34519) begin
		isPrime = 1;
	end	else if (num==16'd34537) begin
		isPrime = 1;
	end	else if (num==16'd34543) begin
		isPrime = 1;
	end	else if (num==16'd34549) begin
		isPrime = 1;
	end	else if (num==16'd34583) begin
		isPrime = 1;
	end	else if (num==16'd34589) begin
		isPrime = 1;
	end	else if (num==16'd34591) begin
		isPrime = 1;
	end	else if (num==16'd34603) begin
		isPrime = 1;
	end	else if (num==16'd34607) begin
		isPrime = 1;
	end	else if (num==16'd34613) begin
		isPrime = 1;
	end	else if (num==16'd34631) begin
		isPrime = 1;
	end	else if (num==16'd34649) begin
		isPrime = 1;
	end	else if (num==16'd34651) begin
		isPrime = 1;
	end	else if (num==16'd34667) begin
		isPrime = 1;
	end	else if (num==16'd34673) begin
		isPrime = 1;
	end	else if (num==16'd34679) begin
		isPrime = 1;
	end	else if (num==16'd34687) begin
		isPrime = 1;
	end	else if (num==16'd34693) begin
		isPrime = 1;
	end	else if (num==16'd34703) begin
		isPrime = 1;
	end	else if (num==16'd34721) begin
		isPrime = 1;
	end	else if (num==16'd34729) begin
		isPrime = 1;
	end	else if (num==16'd34739) begin
		isPrime = 1;
	end	else if (num==16'd34747) begin
		isPrime = 1;
	end	else if (num==16'd34757) begin
		isPrime = 1;
	end	else if (num==16'd34759) begin
		isPrime = 1;
	end	else if (num==16'd34763) begin
		isPrime = 1;
	end	else if (num==16'd34781) begin
		isPrime = 1;
	end	else if (num==16'd34807) begin
		isPrime = 1;
	end	else if (num==16'd34819) begin
		isPrime = 1;
	end	else if (num==16'd34841) begin
		isPrime = 1;
	end	else if (num==16'd34843) begin
		isPrime = 1;
	end	else if (num==16'd34847) begin
		isPrime = 1;
	end	else if (num==16'd34849) begin
		isPrime = 1;
	end	else if (num==16'd34871) begin
		isPrime = 1;
	end	else if (num==16'd34877) begin
		isPrime = 1;
	end	else if (num==16'd34883) begin
		isPrime = 1;
	end	else if (num==16'd34897) begin
		isPrime = 1;
	end	else if (num==16'd34913) begin
		isPrime = 1;
	end	else if (num==16'd34919) begin
		isPrime = 1;
	end	else if (num==16'd34939) begin
		isPrime = 1;
	end	else if (num==16'd34949) begin
		isPrime = 1;
	end	else if (num==16'd34961) begin
		isPrime = 1;
	end	else if (num==16'd34963) begin
		isPrime = 1;
	end	else if (num==16'd34981) begin
		isPrime = 1;
	end	else if (num==16'd35023) begin
		isPrime = 1;
	end	else if (num==16'd35027) begin
		isPrime = 1;
	end	else if (num==16'd35051) begin
		isPrime = 1;
	end	else if (num==16'd35053) begin
		isPrime = 1;
	end	else if (num==16'd35059) begin
		isPrime = 1;
	end	else if (num==16'd35069) begin
		isPrime = 1;
	end	else if (num==16'd35081) begin
		isPrime = 1;
	end	else if (num==16'd35083) begin
		isPrime = 1;
	end	else if (num==16'd35089) begin
		isPrime = 1;
	end	else if (num==16'd35099) begin
		isPrime = 1;
	end	else if (num==16'd35107) begin
		isPrime = 1;
	end	else if (num==16'd35111) begin
		isPrime = 1;
	end	else if (num==16'd35117) begin
		isPrime = 1;
	end	else if (num==16'd35129) begin
		isPrime = 1;
	end	else if (num==16'd35141) begin
		isPrime = 1;
	end	else if (num==16'd35149) begin
		isPrime = 1;
	end	else if (num==16'd35153) begin
		isPrime = 1;
	end	else if (num==16'd35159) begin
		isPrime = 1;
	end	else if (num==16'd35171) begin
		isPrime = 1;
	end	else if (num==16'd35201) begin
		isPrime = 1;
	end	else if (num==16'd35221) begin
		isPrime = 1;
	end	else if (num==16'd35227) begin
		isPrime = 1;
	end	else if (num==16'd35251) begin
		isPrime = 1;
	end	else if (num==16'd35257) begin
		isPrime = 1;
	end	else if (num==16'd35267) begin
		isPrime = 1;
	end	else if (num==16'd35279) begin
		isPrime = 1;
	end	else if (num==16'd35281) begin
		isPrime = 1;
	end	else if (num==16'd35291) begin
		isPrime = 1;
	end	else if (num==16'd35311) begin
		isPrime = 1;
	end	else if (num==16'd35317) begin
		isPrime = 1;
	end	else if (num==16'd35323) begin
		isPrime = 1;
	end	else if (num==16'd35327) begin
		isPrime = 1;
	end	else if (num==16'd35339) begin
		isPrime = 1;
	end	else if (num==16'd35353) begin
		isPrime = 1;
	end	else if (num==16'd35363) begin
		isPrime = 1;
	end	else if (num==16'd35381) begin
		isPrime = 1;
	end	else if (num==16'd35393) begin
		isPrime = 1;
	end	else if (num==16'd35401) begin
		isPrime = 1;
	end	else if (num==16'd35407) begin
		isPrime = 1;
	end	else if (num==16'd35419) begin
		isPrime = 1;
	end	else if (num==16'd35423) begin
		isPrime = 1;
	end	else if (num==16'd35437) begin
		isPrime = 1;
	end	else if (num==16'd35447) begin
		isPrime = 1;
	end	else if (num==16'd35449) begin
		isPrime = 1;
	end	else if (num==16'd35461) begin
		isPrime = 1;
	end	else if (num==16'd35491) begin
		isPrime = 1;
	end	else if (num==16'd35507) begin
		isPrime = 1;
	end	else if (num==16'd35509) begin
		isPrime = 1;
	end	else if (num==16'd35521) begin
		isPrime = 1;
	end	else if (num==16'd35527) begin
		isPrime = 1;
	end	else if (num==16'd35531) begin
		isPrime = 1;
	end	else if (num==16'd35533) begin
		isPrime = 1;
	end	else if (num==16'd35537) begin
		isPrime = 1;
	end	else if (num==16'd35543) begin
		isPrime = 1;
	end	else if (num==16'd35569) begin
		isPrime = 1;
	end	else if (num==16'd35573) begin
		isPrime = 1;
	end	else if (num==16'd35591) begin
		isPrime = 1;
	end	else if (num==16'd35593) begin
		isPrime = 1;
	end	else if (num==16'd35597) begin
		isPrime = 1;
	end	else if (num==16'd35603) begin
		isPrime = 1;
	end	else if (num==16'd35617) begin
		isPrime = 1;
	end	else if (num==16'd35671) begin
		isPrime = 1;
	end	else if (num==16'd35677) begin
		isPrime = 1;
	end	else if (num==16'd35729) begin
		isPrime = 1;
	end	else if (num==16'd35731) begin
		isPrime = 1;
	end	else if (num==16'd35747) begin
		isPrime = 1;
	end	else if (num==16'd35753) begin
		isPrime = 1;
	end	else if (num==16'd35759) begin
		isPrime = 1;
	end	else if (num==16'd35771) begin
		isPrime = 1;
	end	else if (num==16'd35797) begin
		isPrime = 1;
	end	else if (num==16'd35801) begin
		isPrime = 1;
	end	else if (num==16'd35803) begin
		isPrime = 1;
	end	else if (num==16'd35809) begin
		isPrime = 1;
	end	else if (num==16'd35831) begin
		isPrime = 1;
	end	else if (num==16'd35837) begin
		isPrime = 1;
	end	else if (num==16'd35839) begin
		isPrime = 1;
	end	else if (num==16'd35851) begin
		isPrime = 1;
	end	else if (num==16'd35863) begin
		isPrime = 1;
	end	else if (num==16'd35869) begin
		isPrime = 1;
	end	else if (num==16'd35879) begin
		isPrime = 1;
	end	else if (num==16'd35897) begin
		isPrime = 1;
	end	else if (num==16'd35899) begin
		isPrime = 1;
	end	else if (num==16'd35911) begin
		isPrime = 1;
	end	else if (num==16'd35923) begin
		isPrime = 1;
	end	else if (num==16'd35933) begin
		isPrime = 1;
	end	else if (num==16'd35951) begin
		isPrime = 1;
	end	else if (num==16'd35963) begin
		isPrime = 1;
	end	else if (num==16'd35969) begin
		isPrime = 1;
	end	else if (num==16'd35977) begin
		isPrime = 1;
	end	else if (num==16'd35983) begin
		isPrime = 1;
	end	else if (num==16'd35993) begin
		isPrime = 1;
	end	else if (num==16'd35999) begin
		isPrime = 1;
	end	else if (num==16'd36007) begin
		isPrime = 1;
	end	else if (num==16'd36011) begin
		isPrime = 1;
	end	else if (num==16'd36013) begin
		isPrime = 1;
	end	else if (num==16'd36017) begin
		isPrime = 1;
	end	else if (num==16'd36037) begin
		isPrime = 1;
	end	else if (num==16'd36061) begin
		isPrime = 1;
	end	else if (num==16'd36067) begin
		isPrime = 1;
	end	else if (num==16'd36073) begin
		isPrime = 1;
	end	else if (num==16'd36083) begin
		isPrime = 1;
	end	else if (num==16'd36097) begin
		isPrime = 1;
	end	else if (num==16'd36107) begin
		isPrime = 1;
	end	else if (num==16'd36109) begin
		isPrime = 1;
	end	else if (num==16'd36131) begin
		isPrime = 1;
	end	else if (num==16'd36137) begin
		isPrime = 1;
	end	else if (num==16'd36151) begin
		isPrime = 1;
	end	else if (num==16'd36161) begin
		isPrime = 1;
	end	else if (num==16'd36187) begin
		isPrime = 1;
	end	else if (num==16'd36191) begin
		isPrime = 1;
	end	else if (num==16'd36209) begin
		isPrime = 1;
	end	else if (num==16'd36217) begin
		isPrime = 1;
	end	else if (num==16'd36229) begin
		isPrime = 1;
	end	else if (num==16'd36241) begin
		isPrime = 1;
	end	else if (num==16'd36251) begin
		isPrime = 1;
	end	else if (num==16'd36263) begin
		isPrime = 1;
	end	else if (num==16'd36269) begin
		isPrime = 1;
	end	else if (num==16'd36277) begin
		isPrime = 1;
	end	else if (num==16'd36293) begin
		isPrime = 1;
	end	else if (num==16'd36299) begin
		isPrime = 1;
	end	else if (num==16'd36307) begin
		isPrime = 1;
	end	else if (num==16'd36313) begin
		isPrime = 1;
	end	else if (num==16'd36319) begin
		isPrime = 1;
	end	else if (num==16'd36341) begin
		isPrime = 1;
	end	else if (num==16'd36343) begin
		isPrime = 1;
	end	else if (num==16'd36353) begin
		isPrime = 1;
	end	else if (num==16'd36373) begin
		isPrime = 1;
	end	else if (num==16'd36383) begin
		isPrime = 1;
	end	else if (num==16'd36389) begin
		isPrime = 1;
	end	else if (num==16'd36433) begin
		isPrime = 1;
	end	else if (num==16'd36451) begin
		isPrime = 1;
	end	else if (num==16'd36457) begin
		isPrime = 1;
	end	else if (num==16'd36467) begin
		isPrime = 1;
	end	else if (num==16'd36469) begin
		isPrime = 1;
	end	else if (num==16'd36473) begin
		isPrime = 1;
	end	else if (num==16'd36479) begin
		isPrime = 1;
	end	else if (num==16'd36493) begin
		isPrime = 1;
	end	else if (num==16'd36497) begin
		isPrime = 1;
	end	else if (num==16'd36523) begin
		isPrime = 1;
	end	else if (num==16'd36527) begin
		isPrime = 1;
	end	else if (num==16'd36529) begin
		isPrime = 1;
	end	else if (num==16'd36541) begin
		isPrime = 1;
	end	else if (num==16'd36551) begin
		isPrime = 1;
	end	else if (num==16'd36559) begin
		isPrime = 1;
	end	else if (num==16'd36563) begin
		isPrime = 1;
	end	else if (num==16'd36571) begin
		isPrime = 1;
	end	else if (num==16'd36583) begin
		isPrime = 1;
	end	else if (num==16'd36587) begin
		isPrime = 1;
	end	else if (num==16'd36599) begin
		isPrime = 1;
	end	else if (num==16'd36607) begin
		isPrime = 1;
	end	else if (num==16'd36629) begin
		isPrime = 1;
	end	else if (num==16'd36637) begin
		isPrime = 1;
	end	else if (num==16'd36643) begin
		isPrime = 1;
	end	else if (num==16'd36653) begin
		isPrime = 1;
	end	else if (num==16'd36671) begin
		isPrime = 1;
	end	else if (num==16'd36677) begin
		isPrime = 1;
	end	else if (num==16'd36683) begin
		isPrime = 1;
	end	else if (num==16'd36691) begin
		isPrime = 1;
	end	else if (num==16'd36697) begin
		isPrime = 1;
	end	else if (num==16'd36709) begin
		isPrime = 1;
	end	else if (num==16'd36713) begin
		isPrime = 1;
	end	else if (num==16'd36721) begin
		isPrime = 1;
	end	else if (num==16'd36739) begin
		isPrime = 1;
	end	else if (num==16'd36749) begin
		isPrime = 1;
	end	else if (num==16'd36761) begin
		isPrime = 1;
	end	else if (num==16'd36767) begin
		isPrime = 1;
	end	else if (num==16'd36779) begin
		isPrime = 1;
	end	else if (num==16'd36781) begin
		isPrime = 1;
	end	else if (num==16'd36787) begin
		isPrime = 1;
	end	else if (num==16'd36791) begin
		isPrime = 1;
	end	else if (num==16'd36793) begin
		isPrime = 1;
	end	else if (num==16'd36809) begin
		isPrime = 1;
	end	else if (num==16'd36821) begin
		isPrime = 1;
	end	else if (num==16'd36833) begin
		isPrime = 1;
	end	else if (num==16'd36847) begin
		isPrime = 1;
	end	else if (num==16'd36857) begin
		isPrime = 1;
	end	else if (num==16'd36871) begin
		isPrime = 1;
	end	else if (num==16'd36877) begin
		isPrime = 1;
	end	else if (num==16'd36887) begin
		isPrime = 1;
	end	else if (num==16'd36899) begin
		isPrime = 1;
	end	else if (num==16'd36901) begin
		isPrime = 1;
	end	else if (num==16'd36913) begin
		isPrime = 1;
	end	else if (num==16'd36919) begin
		isPrime = 1;
	end	else if (num==16'd36923) begin
		isPrime = 1;
	end	else if (num==16'd36929) begin
		isPrime = 1;
	end	else if (num==16'd36931) begin
		isPrime = 1;
	end	else if (num==16'd36943) begin
		isPrime = 1;
	end	else if (num==16'd36947) begin
		isPrime = 1;
	end	else if (num==16'd36973) begin
		isPrime = 1;
	end	else if (num==16'd36979) begin
		isPrime = 1;
	end	else if (num==16'd36997) begin
		isPrime = 1;
	end	else if (num==16'd37003) begin
		isPrime = 1;
	end	else if (num==16'd37013) begin
		isPrime = 1;
	end	else if (num==16'd37019) begin
		isPrime = 1;
	end	else if (num==16'd37021) begin
		isPrime = 1;
	end	else if (num==16'd37039) begin
		isPrime = 1;
	end	else if (num==16'd37049) begin
		isPrime = 1;
	end	else if (num==16'd37057) begin
		isPrime = 1;
	end	else if (num==16'd37061) begin
		isPrime = 1;
	end	else if (num==16'd37087) begin
		isPrime = 1;
	end	else if (num==16'd37097) begin
		isPrime = 1;
	end	else if (num==16'd37117) begin
		isPrime = 1;
	end	else if (num==16'd37123) begin
		isPrime = 1;
	end	else if (num==16'd37139) begin
		isPrime = 1;
	end	else if (num==16'd37159) begin
		isPrime = 1;
	end	else if (num==16'd37171) begin
		isPrime = 1;
	end	else if (num==16'd37181) begin
		isPrime = 1;
	end	else if (num==16'd37189) begin
		isPrime = 1;
	end	else if (num==16'd37199) begin
		isPrime = 1;
	end	else if (num==16'd37201) begin
		isPrime = 1;
	end	else if (num==16'd37217) begin
		isPrime = 1;
	end	else if (num==16'd37223) begin
		isPrime = 1;
	end	else if (num==16'd37243) begin
		isPrime = 1;
	end	else if (num==16'd37253) begin
		isPrime = 1;
	end	else if (num==16'd37273) begin
		isPrime = 1;
	end	else if (num==16'd37277) begin
		isPrime = 1;
	end	else if (num==16'd37307) begin
		isPrime = 1;
	end	else if (num==16'd37309) begin
		isPrime = 1;
	end	else if (num==16'd37313) begin
		isPrime = 1;
	end	else if (num==16'd37321) begin
		isPrime = 1;
	end	else if (num==16'd37337) begin
		isPrime = 1;
	end	else if (num==16'd37339) begin
		isPrime = 1;
	end	else if (num==16'd37357) begin
		isPrime = 1;
	end	else if (num==16'd37361) begin
		isPrime = 1;
	end	else if (num==16'd37363) begin
		isPrime = 1;
	end	else if (num==16'd37369) begin
		isPrime = 1;
	end	else if (num==16'd37379) begin
		isPrime = 1;
	end	else if (num==16'd37397) begin
		isPrime = 1;
	end	else if (num==16'd37409) begin
		isPrime = 1;
	end	else if (num==16'd37423) begin
		isPrime = 1;
	end	else if (num==16'd37441) begin
		isPrime = 1;
	end	else if (num==16'd37447) begin
		isPrime = 1;
	end	else if (num==16'd37463) begin
		isPrime = 1;
	end	else if (num==16'd37483) begin
		isPrime = 1;
	end	else if (num==16'd37489) begin
		isPrime = 1;
	end	else if (num==16'd37493) begin
		isPrime = 1;
	end	else if (num==16'd37501) begin
		isPrime = 1;
	end	else if (num==16'd37507) begin
		isPrime = 1;
	end	else if (num==16'd37511) begin
		isPrime = 1;
	end	else if (num==16'd37517) begin
		isPrime = 1;
	end	else if (num==16'd37529) begin
		isPrime = 1;
	end	else if (num==16'd37537) begin
		isPrime = 1;
	end	else if (num==16'd37547) begin
		isPrime = 1;
	end	else if (num==16'd37549) begin
		isPrime = 1;
	end	else if (num==16'd37561) begin
		isPrime = 1;
	end	else if (num==16'd37567) begin
		isPrime = 1;
	end	else if (num==16'd37571) begin
		isPrime = 1;
	end	else if (num==16'd37573) begin
		isPrime = 1;
	end	else if (num==16'd37579) begin
		isPrime = 1;
	end	else if (num==16'd37589) begin
		isPrime = 1;
	end	else if (num==16'd37591) begin
		isPrime = 1;
	end	else if (num==16'd37607) begin
		isPrime = 1;
	end	else if (num==16'd37619) begin
		isPrime = 1;
	end	else if (num==16'd37633) begin
		isPrime = 1;
	end	else if (num==16'd37643) begin
		isPrime = 1;
	end	else if (num==16'd37649) begin
		isPrime = 1;
	end	else if (num==16'd37657) begin
		isPrime = 1;
	end	else if (num==16'd37663) begin
		isPrime = 1;
	end	else if (num==16'd37691) begin
		isPrime = 1;
	end	else if (num==16'd37693) begin
		isPrime = 1;
	end	else if (num==16'd37699) begin
		isPrime = 1;
	end	else if (num==16'd37717) begin
		isPrime = 1;
	end	else if (num==16'd37747) begin
		isPrime = 1;
	end	else if (num==16'd37781) begin
		isPrime = 1;
	end	else if (num==16'd37783) begin
		isPrime = 1;
	end	else if (num==16'd37799) begin
		isPrime = 1;
	end	else if (num==16'd37811) begin
		isPrime = 1;
	end	else if (num==16'd37813) begin
		isPrime = 1;
	end	else if (num==16'd37831) begin
		isPrime = 1;
	end	else if (num==16'd37847) begin
		isPrime = 1;
	end	else if (num==16'd37853) begin
		isPrime = 1;
	end	else if (num==16'd37861) begin
		isPrime = 1;
	end	else if (num==16'd37871) begin
		isPrime = 1;
	end	else if (num==16'd37879) begin
		isPrime = 1;
	end	else if (num==16'd37889) begin
		isPrime = 1;
	end	else if (num==16'd37897) begin
		isPrime = 1;
	end	else if (num==16'd37907) begin
		isPrime = 1;
	end	else if (num==16'd37951) begin
		isPrime = 1;
	end	else if (num==16'd37957) begin
		isPrime = 1;
	end	else if (num==16'd37963) begin
		isPrime = 1;
	end	else if (num==16'd37967) begin
		isPrime = 1;
	end	else if (num==16'd37987) begin
		isPrime = 1;
	end	else if (num==16'd37991) begin
		isPrime = 1;
	end	else if (num==16'd37993) begin
		isPrime = 1;
	end	else if (num==16'd37997) begin
		isPrime = 1;
	end	else if (num==16'd38011) begin
		isPrime = 1;
	end	else if (num==16'd38039) begin
		isPrime = 1;
	end	else if (num==16'd38047) begin
		isPrime = 1;
	end	else if (num==16'd38053) begin
		isPrime = 1;
	end	else if (num==16'd38069) begin
		isPrime = 1;
	end	else if (num==16'd38083) begin
		isPrime = 1;
	end	else if (num==16'd38113) begin
		isPrime = 1;
	end	else if (num==16'd38119) begin
		isPrime = 1;
	end	else if (num==16'd38149) begin
		isPrime = 1;
	end	else if (num==16'd38153) begin
		isPrime = 1;
	end	else if (num==16'd38167) begin
		isPrime = 1;
	end	else if (num==16'd38177) begin
		isPrime = 1;
	end	else if (num==16'd38183) begin
		isPrime = 1;
	end	else if (num==16'd38189) begin
		isPrime = 1;
	end	else if (num==16'd38197) begin
		isPrime = 1;
	end	else if (num==16'd38201) begin
		isPrime = 1;
	end	else if (num==16'd38219) begin
		isPrime = 1;
	end	else if (num==16'd38231) begin
		isPrime = 1;
	end	else if (num==16'd38237) begin
		isPrime = 1;
	end	else if (num==16'd38239) begin
		isPrime = 1;
	end	else if (num==16'd38261) begin
		isPrime = 1;
	end	else if (num==16'd38273) begin
		isPrime = 1;
	end	else if (num==16'd38281) begin
		isPrime = 1;
	end	else if (num==16'd38287) begin
		isPrime = 1;
	end	else if (num==16'd38299) begin
		isPrime = 1;
	end	else if (num==16'd38303) begin
		isPrime = 1;
	end	else if (num==16'd38317) begin
		isPrime = 1;
	end	else if (num==16'd38321) begin
		isPrime = 1;
	end	else if (num==16'd38327) begin
		isPrime = 1;
	end	else if (num==16'd38329) begin
		isPrime = 1;
	end	else if (num==16'd38333) begin
		isPrime = 1;
	end	else if (num==16'd38351) begin
		isPrime = 1;
	end	else if (num==16'd38371) begin
		isPrime = 1;
	end	else if (num==16'd38377) begin
		isPrime = 1;
	end	else if (num==16'd38393) begin
		isPrime = 1;
	end	else if (num==16'd38431) begin
		isPrime = 1;
	end	else if (num==16'd38447) begin
		isPrime = 1;
	end	else if (num==16'd38449) begin
		isPrime = 1;
	end	else if (num==16'd38453) begin
		isPrime = 1;
	end	else if (num==16'd38459) begin
		isPrime = 1;
	end	else if (num==16'd38461) begin
		isPrime = 1;
	end	else if (num==16'd38501) begin
		isPrime = 1;
	end	else if (num==16'd38543) begin
		isPrime = 1;
	end	else if (num==16'd38557) begin
		isPrime = 1;
	end	else if (num==16'd38561) begin
		isPrime = 1;
	end	else if (num==16'd38567) begin
		isPrime = 1;
	end	else if (num==16'd38569) begin
		isPrime = 1;
	end	else if (num==16'd38593) begin
		isPrime = 1;
	end	else if (num==16'd38603) begin
		isPrime = 1;
	end	else if (num==16'd38609) begin
		isPrime = 1;
	end	else if (num==16'd38611) begin
		isPrime = 1;
	end	else if (num==16'd38629) begin
		isPrime = 1;
	end	else if (num==16'd38639) begin
		isPrime = 1;
	end	else if (num==16'd38651) begin
		isPrime = 1;
	end	else if (num==16'd38653) begin
		isPrime = 1;
	end	else if (num==16'd38669) begin
		isPrime = 1;
	end	else if (num==16'd38671) begin
		isPrime = 1;
	end	else if (num==16'd38677) begin
		isPrime = 1;
	end	else if (num==16'd38693) begin
		isPrime = 1;
	end	else if (num==16'd38699) begin
		isPrime = 1;
	end	else if (num==16'd38707) begin
		isPrime = 1;
	end	else if (num==16'd38711) begin
		isPrime = 1;
	end	else if (num==16'd38713) begin
		isPrime = 1;
	end	else if (num==16'd38723) begin
		isPrime = 1;
	end	else if (num==16'd38729) begin
		isPrime = 1;
	end	else if (num==16'd38737) begin
		isPrime = 1;
	end	else if (num==16'd38747) begin
		isPrime = 1;
	end	else if (num==16'd38749) begin
		isPrime = 1;
	end	else if (num==16'd38767) begin
		isPrime = 1;
	end	else if (num==16'd38783) begin
		isPrime = 1;
	end	else if (num==16'd38791) begin
		isPrime = 1;
	end	else if (num==16'd38803) begin
		isPrime = 1;
	end	else if (num==16'd38821) begin
		isPrime = 1;
	end	else if (num==16'd38833) begin
		isPrime = 1;
	end	else if (num==16'd38839) begin
		isPrime = 1;
	end	else if (num==16'd38851) begin
		isPrime = 1;
	end	else if (num==16'd38861) begin
		isPrime = 1;
	end	else if (num==16'd38867) begin
		isPrime = 1;
	end	else if (num==16'd38873) begin
		isPrime = 1;
	end	else if (num==16'd38891) begin
		isPrime = 1;
	end	else if (num==16'd38903) begin
		isPrime = 1;
	end	else if (num==16'd38917) begin
		isPrime = 1;
	end	else if (num==16'd38921) begin
		isPrime = 1;
	end	else if (num==16'd38923) begin
		isPrime = 1;
	end	else if (num==16'd38933) begin
		isPrime = 1;
	end	else if (num==16'd38953) begin
		isPrime = 1;
	end	else if (num==16'd38959) begin
		isPrime = 1;
	end	else if (num==16'd38971) begin
		isPrime = 1;
	end	else if (num==16'd38977) begin
		isPrime = 1;
	end	else if (num==16'd38993) begin
		isPrime = 1;
	end	else if (num==16'd39019) begin
		isPrime = 1;
	end	else if (num==16'd39023) begin
		isPrime = 1;
	end	else if (num==16'd39041) begin
		isPrime = 1;
	end	else if (num==16'd39043) begin
		isPrime = 1;
	end	else if (num==16'd39047) begin
		isPrime = 1;
	end	else if (num==16'd39079) begin
		isPrime = 1;
	end	else if (num==16'd39089) begin
		isPrime = 1;
	end	else if (num==16'd39097) begin
		isPrime = 1;
	end	else if (num==16'd39103) begin
		isPrime = 1;
	end	else if (num==16'd39107) begin
		isPrime = 1;
	end	else if (num==16'd39113) begin
		isPrime = 1;
	end	else if (num==16'd39119) begin
		isPrime = 1;
	end	else if (num==16'd39133) begin
		isPrime = 1;
	end	else if (num==16'd39139) begin
		isPrime = 1;
	end	else if (num==16'd39157) begin
		isPrime = 1;
	end	else if (num==16'd39161) begin
		isPrime = 1;
	end	else if (num==16'd39163) begin
		isPrime = 1;
	end	else if (num==16'd39181) begin
		isPrime = 1;
	end	else if (num==16'd39191) begin
		isPrime = 1;
	end	else if (num==16'd39199) begin
		isPrime = 1;
	end	else if (num==16'd39209) begin
		isPrime = 1;
	end	else if (num==16'd39217) begin
		isPrime = 1;
	end	else if (num==16'd39227) begin
		isPrime = 1;
	end	else if (num==16'd39229) begin
		isPrime = 1;
	end	else if (num==16'd39233) begin
		isPrime = 1;
	end	else if (num==16'd39239) begin
		isPrime = 1;
	end	else if (num==16'd39241) begin
		isPrime = 1;
	end	else if (num==16'd39251) begin
		isPrime = 1;
	end	else if (num==16'd39293) begin
		isPrime = 1;
	end	else if (num==16'd39301) begin
		isPrime = 1;
	end	else if (num==16'd39313) begin
		isPrime = 1;
	end	else if (num==16'd39317) begin
		isPrime = 1;
	end	else if (num==16'd39323) begin
		isPrime = 1;
	end	else if (num==16'd39341) begin
		isPrime = 1;
	end	else if (num==16'd39343) begin
		isPrime = 1;
	end	else if (num==16'd39359) begin
		isPrime = 1;
	end	else if (num==16'd39367) begin
		isPrime = 1;
	end	else if (num==16'd39371) begin
		isPrime = 1;
	end	else if (num==16'd39373) begin
		isPrime = 1;
	end	else if (num==16'd39383) begin
		isPrime = 1;
	end	else if (num==16'd39397) begin
		isPrime = 1;
	end	else if (num==16'd39409) begin
		isPrime = 1;
	end	else if (num==16'd39419) begin
		isPrime = 1;
	end	else if (num==16'd39439) begin
		isPrime = 1;
	end	else if (num==16'd39443) begin
		isPrime = 1;
	end	else if (num==16'd39451) begin
		isPrime = 1;
	end	else if (num==16'd39461) begin
		isPrime = 1;
	end	else if (num==16'd39499) begin
		isPrime = 1;
	end	else if (num==16'd39503) begin
		isPrime = 1;
	end	else if (num==16'd39509) begin
		isPrime = 1;
	end	else if (num==16'd39511) begin
		isPrime = 1;
	end	else if (num==16'd39521) begin
		isPrime = 1;
	end	else if (num==16'd39541) begin
		isPrime = 1;
	end	else if (num==16'd39551) begin
		isPrime = 1;
	end	else if (num==16'd39563) begin
		isPrime = 1;
	end	else if (num==16'd39569) begin
		isPrime = 1;
	end	else if (num==16'd39581) begin
		isPrime = 1;
	end	else if (num==16'd39607) begin
		isPrime = 1;
	end	else if (num==16'd39619) begin
		isPrime = 1;
	end	else if (num==16'd39623) begin
		isPrime = 1;
	end	else if (num==16'd39631) begin
		isPrime = 1;
	end	else if (num==16'd39659) begin
		isPrime = 1;
	end	else if (num==16'd39667) begin
		isPrime = 1;
	end	else if (num==16'd39671) begin
		isPrime = 1;
	end	else if (num==16'd39679) begin
		isPrime = 1;
	end	else if (num==16'd39703) begin
		isPrime = 1;
	end	else if (num==16'd39709) begin
		isPrime = 1;
	end	else if (num==16'd39719) begin
		isPrime = 1;
	end	else if (num==16'd39727) begin
		isPrime = 1;
	end	else if (num==16'd39733) begin
		isPrime = 1;
	end	else if (num==16'd39749) begin
		isPrime = 1;
	end	else if (num==16'd39761) begin
		isPrime = 1;
	end	else if (num==16'd39769) begin
		isPrime = 1;
	end	else if (num==16'd39779) begin
		isPrime = 1;
	end	else if (num==16'd39791) begin
		isPrime = 1;
	end	else if (num==16'd39799) begin
		isPrime = 1;
	end	else if (num==16'd39821) begin
		isPrime = 1;
	end	else if (num==16'd39827) begin
		isPrime = 1;
	end	else if (num==16'd39829) begin
		isPrime = 1;
	end	else if (num==16'd39839) begin
		isPrime = 1;
	end	else if (num==16'd39841) begin
		isPrime = 1;
	end	else if (num==16'd39847) begin
		isPrime = 1;
	end	else if (num==16'd39857) begin
		isPrime = 1;
	end	else if (num==16'd39863) begin
		isPrime = 1;
	end	else if (num==16'd39869) begin
		isPrime = 1;
	end	else if (num==16'd39877) begin
		isPrime = 1;
	end	else if (num==16'd39883) begin
		isPrime = 1;
	end	else if (num==16'd39887) begin
		isPrime = 1;
	end	else if (num==16'd39901) begin
		isPrime = 1;
	end	else if (num==16'd39929) begin
		isPrime = 1;
	end	else if (num==16'd39937) begin
		isPrime = 1;
	end	else if (num==16'd39953) begin
		isPrime = 1;
	end	else if (num==16'd39971) begin
		isPrime = 1;
	end	else if (num==16'd39979) begin
		isPrime = 1;
	end	else if (num==16'd39983) begin
		isPrime = 1;
	end	else if (num==16'd39989) begin
		isPrime = 1;
	end	else if (num==16'd40009) begin
		isPrime = 1;
	end	else if (num==16'd40013) begin
		isPrime = 1;
	end	else if (num==16'd40031) begin
		isPrime = 1;
	end	else if (num==16'd40037) begin
		isPrime = 1;
	end	else if (num==16'd40039) begin
		isPrime = 1;
	end	else if (num==16'd40063) begin
		isPrime = 1;
	end	else if (num==16'd40087) begin
		isPrime = 1;
	end	else if (num==16'd40093) begin
		isPrime = 1;
	end	else if (num==16'd40099) begin
		isPrime = 1;
	end	else if (num==16'd40111) begin
		isPrime = 1;
	end	else if (num==16'd40123) begin
		isPrime = 1;
	end	else if (num==16'd40127) begin
		isPrime = 1;
	end	else if (num==16'd40129) begin
		isPrime = 1;
	end	else if (num==16'd40151) begin
		isPrime = 1;
	end	else if (num==16'd40153) begin
		isPrime = 1;
	end	else if (num==16'd40163) begin
		isPrime = 1;
	end	else if (num==16'd40169) begin
		isPrime = 1;
	end	else if (num==16'd40177) begin
		isPrime = 1;
	end	else if (num==16'd40189) begin
		isPrime = 1;
	end	else if (num==16'd40193) begin
		isPrime = 1;
	end	else if (num==16'd40213) begin
		isPrime = 1;
	end	else if (num==16'd40231) begin
		isPrime = 1;
	end	else if (num==16'd40237) begin
		isPrime = 1;
	end	else if (num==16'd40241) begin
		isPrime = 1;
	end	else if (num==16'd40253) begin
		isPrime = 1;
	end	else if (num==16'd40277) begin
		isPrime = 1;
	end	else if (num==16'd40283) begin
		isPrime = 1;
	end	else if (num==16'd40289) begin
		isPrime = 1;
	end	else if (num==16'd40343) begin
		isPrime = 1;
	end	else if (num==16'd40351) begin
		isPrime = 1;
	end	else if (num==16'd40357) begin
		isPrime = 1;
	end	else if (num==16'd40361) begin
		isPrime = 1;
	end	else if (num==16'd40387) begin
		isPrime = 1;
	end	else if (num==16'd40423) begin
		isPrime = 1;
	end	else if (num==16'd40427) begin
		isPrime = 1;
	end	else if (num==16'd40429) begin
		isPrime = 1;
	end	else if (num==16'd40433) begin
		isPrime = 1;
	end	else if (num==16'd40459) begin
		isPrime = 1;
	end	else if (num==16'd40471) begin
		isPrime = 1;
	end	else if (num==16'd40483) begin
		isPrime = 1;
	end	else if (num==16'd40487) begin
		isPrime = 1;
	end	else if (num==16'd40493) begin
		isPrime = 1;
	end	else if (num==16'd40499) begin
		isPrime = 1;
	end	else if (num==16'd40507) begin
		isPrime = 1;
	end	else if (num==16'd40519) begin
		isPrime = 1;
	end	else if (num==16'd40529) begin
		isPrime = 1;
	end	else if (num==16'd40531) begin
		isPrime = 1;
	end	else if (num==16'd40543) begin
		isPrime = 1;
	end	else if (num==16'd40559) begin
		isPrime = 1;
	end	else if (num==16'd40577) begin
		isPrime = 1;
	end	else if (num==16'd40583) begin
		isPrime = 1;
	end	else if (num==16'd40591) begin
		isPrime = 1;
	end	else if (num==16'd40597) begin
		isPrime = 1;
	end	else if (num==16'd40609) begin
		isPrime = 1;
	end	else if (num==16'd40627) begin
		isPrime = 1;
	end	else if (num==16'd40637) begin
		isPrime = 1;
	end	else if (num==16'd40639) begin
		isPrime = 1;
	end	else if (num==16'd40693) begin
		isPrime = 1;
	end	else if (num==16'd40697) begin
		isPrime = 1;
	end	else if (num==16'd40699) begin
		isPrime = 1;
	end	else if (num==16'd40709) begin
		isPrime = 1;
	end	else if (num==16'd40739) begin
		isPrime = 1;
	end	else if (num==16'd40751) begin
		isPrime = 1;
	end	else if (num==16'd40759) begin
		isPrime = 1;
	end	else if (num==16'd40763) begin
		isPrime = 1;
	end	else if (num==16'd40771) begin
		isPrime = 1;
	end	else if (num==16'd40787) begin
		isPrime = 1;
	end	else if (num==16'd40801) begin
		isPrime = 1;
	end	else if (num==16'd40813) begin
		isPrime = 1;
	end	else if (num==16'd40819) begin
		isPrime = 1;
	end	else if (num==16'd40823) begin
		isPrime = 1;
	end	else if (num==16'd40829) begin
		isPrime = 1;
	end	else if (num==16'd40841) begin
		isPrime = 1;
	end	else if (num==16'd40847) begin
		isPrime = 1;
	end	else if (num==16'd40849) begin
		isPrime = 1;
	end	else if (num==16'd40853) begin
		isPrime = 1;
	end	else if (num==16'd40867) begin
		isPrime = 1;
	end	else if (num==16'd40879) begin
		isPrime = 1;
	end	else if (num==16'd40883) begin
		isPrime = 1;
	end	else if (num==16'd40897) begin
		isPrime = 1;
	end	else if (num==16'd40903) begin
		isPrime = 1;
	end	else if (num==16'd40927) begin
		isPrime = 1;
	end	else if (num==16'd40933) begin
		isPrime = 1;
	end	else if (num==16'd40939) begin
		isPrime = 1;
	end	else if (num==16'd40949) begin
		isPrime = 1;
	end	else if (num==16'd40961) begin
		isPrime = 1;
	end	else if (num==16'd40973) begin
		isPrime = 1;
	end	else if (num==16'd40993) begin
		isPrime = 1;
	end	else if (num==16'd41011) begin
		isPrime = 1;
	end	else if (num==16'd41017) begin
		isPrime = 1;
	end	else if (num==16'd41023) begin
		isPrime = 1;
	end	else if (num==16'd41039) begin
		isPrime = 1;
	end	else if (num==16'd41047) begin
		isPrime = 1;
	end	else if (num==16'd41051) begin
		isPrime = 1;
	end	else if (num==16'd41057) begin
		isPrime = 1;
	end	else if (num==16'd41077) begin
		isPrime = 1;
	end	else if (num==16'd41081) begin
		isPrime = 1;
	end	else if (num==16'd41113) begin
		isPrime = 1;
	end	else if (num==16'd41117) begin
		isPrime = 1;
	end	else if (num==16'd41131) begin
		isPrime = 1;
	end	else if (num==16'd41141) begin
		isPrime = 1;
	end	else if (num==16'd41143) begin
		isPrime = 1;
	end	else if (num==16'd41149) begin
		isPrime = 1;
	end	else if (num==16'd41161) begin
		isPrime = 1;
	end	else if (num==16'd41177) begin
		isPrime = 1;
	end	else if (num==16'd41179) begin
		isPrime = 1;
	end	else if (num==16'd41183) begin
		isPrime = 1;
	end	else if (num==16'd41189) begin
		isPrime = 1;
	end	else if (num==16'd41201) begin
		isPrime = 1;
	end	else if (num==16'd41203) begin
		isPrime = 1;
	end	else if (num==16'd41213) begin
		isPrime = 1;
	end	else if (num==16'd41221) begin
		isPrime = 1;
	end	else if (num==16'd41227) begin
		isPrime = 1;
	end	else if (num==16'd41231) begin
		isPrime = 1;
	end	else if (num==16'd41233) begin
		isPrime = 1;
	end	else if (num==16'd41243) begin
		isPrime = 1;
	end	else if (num==16'd41257) begin
		isPrime = 1;
	end	else if (num==16'd41263) begin
		isPrime = 1;
	end	else if (num==16'd41269) begin
		isPrime = 1;
	end	else if (num==16'd41281) begin
		isPrime = 1;
	end	else if (num==16'd41299) begin
		isPrime = 1;
	end	else if (num==16'd41333) begin
		isPrime = 1;
	end	else if (num==16'd41341) begin
		isPrime = 1;
	end	else if (num==16'd41351) begin
		isPrime = 1;
	end	else if (num==16'd41357) begin
		isPrime = 1;
	end	else if (num==16'd41381) begin
		isPrime = 1;
	end	else if (num==16'd41387) begin
		isPrime = 1;
	end	else if (num==16'd41389) begin
		isPrime = 1;
	end	else if (num==16'd41399) begin
		isPrime = 1;
	end	else if (num==16'd41411) begin
		isPrime = 1;
	end	else if (num==16'd41413) begin
		isPrime = 1;
	end	else if (num==16'd41443) begin
		isPrime = 1;
	end	else if (num==16'd41453) begin
		isPrime = 1;
	end	else if (num==16'd41467) begin
		isPrime = 1;
	end	else if (num==16'd41479) begin
		isPrime = 1;
	end	else if (num==16'd41491) begin
		isPrime = 1;
	end	else if (num==16'd41507) begin
		isPrime = 1;
	end	else if (num==16'd41513) begin
		isPrime = 1;
	end	else if (num==16'd41519) begin
		isPrime = 1;
	end	else if (num==16'd41521) begin
		isPrime = 1;
	end	else if (num==16'd41539) begin
		isPrime = 1;
	end	else if (num==16'd41543) begin
		isPrime = 1;
	end	else if (num==16'd41549) begin
		isPrime = 1;
	end	else if (num==16'd41579) begin
		isPrime = 1;
	end	else if (num==16'd41593) begin
		isPrime = 1;
	end	else if (num==16'd41597) begin
		isPrime = 1;
	end	else if (num==16'd41603) begin
		isPrime = 1;
	end	else if (num==16'd41609) begin
		isPrime = 1;
	end	else if (num==16'd41611) begin
		isPrime = 1;
	end	else if (num==16'd41617) begin
		isPrime = 1;
	end	else if (num==16'd41621) begin
		isPrime = 1;
	end	else if (num==16'd41627) begin
		isPrime = 1;
	end	else if (num==16'd41641) begin
		isPrime = 1;
	end	else if (num==16'd41647) begin
		isPrime = 1;
	end	else if (num==16'd41651) begin
		isPrime = 1;
	end	else if (num==16'd41659) begin
		isPrime = 1;
	end	else if (num==16'd41669) begin
		isPrime = 1;
	end	else if (num==16'd41681) begin
		isPrime = 1;
	end	else if (num==16'd41687) begin
		isPrime = 1;
	end	else if (num==16'd41719) begin
		isPrime = 1;
	end	else if (num==16'd41729) begin
		isPrime = 1;
	end	else if (num==16'd41737) begin
		isPrime = 1;
	end	else if (num==16'd41759) begin
		isPrime = 1;
	end	else if (num==16'd41761) begin
		isPrime = 1;
	end	else if (num==16'd41771) begin
		isPrime = 1;
	end	else if (num==16'd41777) begin
		isPrime = 1;
	end	else if (num==16'd41801) begin
		isPrime = 1;
	end	else if (num==16'd41809) begin
		isPrime = 1;
	end	else if (num==16'd41813) begin
		isPrime = 1;
	end	else if (num==16'd41843) begin
		isPrime = 1;
	end	else if (num==16'd41849) begin
		isPrime = 1;
	end	else if (num==16'd41851) begin
		isPrime = 1;
	end	else if (num==16'd41863) begin
		isPrime = 1;
	end	else if (num==16'd41879) begin
		isPrime = 1;
	end	else if (num==16'd41887) begin
		isPrime = 1;
	end	else if (num==16'd41893) begin
		isPrime = 1;
	end	else if (num==16'd41897) begin
		isPrime = 1;
	end	else if (num==16'd41903) begin
		isPrime = 1;
	end	else if (num==16'd41911) begin
		isPrime = 1;
	end	else if (num==16'd41927) begin
		isPrime = 1;
	end	else if (num==16'd41941) begin
		isPrime = 1;
	end	else if (num==16'd41947) begin
		isPrime = 1;
	end	else if (num==16'd41953) begin
		isPrime = 1;
	end	else if (num==16'd41957) begin
		isPrime = 1;
	end	else if (num==16'd41959) begin
		isPrime = 1;
	end	else if (num==16'd41969) begin
		isPrime = 1;
	end	else if (num==16'd41981) begin
		isPrime = 1;
	end	else if (num==16'd41983) begin
		isPrime = 1;
	end	else if (num==16'd41999) begin
		isPrime = 1;
	end	else if (num==16'd42013) begin
		isPrime = 1;
	end	else if (num==16'd42017) begin
		isPrime = 1;
	end	else if (num==16'd42019) begin
		isPrime = 1;
	end	else if (num==16'd42023) begin
		isPrime = 1;
	end	else if (num==16'd42043) begin
		isPrime = 1;
	end	else if (num==16'd42061) begin
		isPrime = 1;
	end	else if (num==16'd42071) begin
		isPrime = 1;
	end	else if (num==16'd42073) begin
		isPrime = 1;
	end	else if (num==16'd42083) begin
		isPrime = 1;
	end	else if (num==16'd42089) begin
		isPrime = 1;
	end	else if (num==16'd42101) begin
		isPrime = 1;
	end	else if (num==16'd42131) begin
		isPrime = 1;
	end	else if (num==16'd42139) begin
		isPrime = 1;
	end	else if (num==16'd42157) begin
		isPrime = 1;
	end	else if (num==16'd42169) begin
		isPrime = 1;
	end	else if (num==16'd42179) begin
		isPrime = 1;
	end	else if (num==16'd42181) begin
		isPrime = 1;
	end	else if (num==16'd42187) begin
		isPrime = 1;
	end	else if (num==16'd42193) begin
		isPrime = 1;
	end	else if (num==16'd42197) begin
		isPrime = 1;
	end	else if (num==16'd42209) begin
		isPrime = 1;
	end	else if (num==16'd42221) begin
		isPrime = 1;
	end	else if (num==16'd42223) begin
		isPrime = 1;
	end	else if (num==16'd42227) begin
		isPrime = 1;
	end	else if (num==16'd42239) begin
		isPrime = 1;
	end	else if (num==16'd42257) begin
		isPrime = 1;
	end	else if (num==16'd42281) begin
		isPrime = 1;
	end	else if (num==16'd42283) begin
		isPrime = 1;
	end	else if (num==16'd42293) begin
		isPrime = 1;
	end	else if (num==16'd42299) begin
		isPrime = 1;
	end	else if (num==16'd42307) begin
		isPrime = 1;
	end	else if (num==16'd42323) begin
		isPrime = 1;
	end	else if (num==16'd42331) begin
		isPrime = 1;
	end	else if (num==16'd42337) begin
		isPrime = 1;
	end	else if (num==16'd42349) begin
		isPrime = 1;
	end	else if (num==16'd42359) begin
		isPrime = 1;
	end	else if (num==16'd42373) begin
		isPrime = 1;
	end	else if (num==16'd42379) begin
		isPrime = 1;
	end	else if (num==16'd42391) begin
		isPrime = 1;
	end	else if (num==16'd42397) begin
		isPrime = 1;
	end	else if (num==16'd42403) begin
		isPrime = 1;
	end	else if (num==16'd42407) begin
		isPrime = 1;
	end	else if (num==16'd42409) begin
		isPrime = 1;
	end	else if (num==16'd42433) begin
		isPrime = 1;
	end	else if (num==16'd42437) begin
		isPrime = 1;
	end	else if (num==16'd42443) begin
		isPrime = 1;
	end	else if (num==16'd42451) begin
		isPrime = 1;
	end	else if (num==16'd42457) begin
		isPrime = 1;
	end	else if (num==16'd42461) begin
		isPrime = 1;
	end	else if (num==16'd42463) begin
		isPrime = 1;
	end	else if (num==16'd42467) begin
		isPrime = 1;
	end	else if (num==16'd42473) begin
		isPrime = 1;
	end	else if (num==16'd42487) begin
		isPrime = 1;
	end	else if (num==16'd42491) begin
		isPrime = 1;
	end	else if (num==16'd42499) begin
		isPrime = 1;
	end	else if (num==16'd42509) begin
		isPrime = 1;
	end	else if (num==16'd42533) begin
		isPrime = 1;
	end	else if (num==16'd42557) begin
		isPrime = 1;
	end	else if (num==16'd42569) begin
		isPrime = 1;
	end	else if (num==16'd42571) begin
		isPrime = 1;
	end	else if (num==16'd42577) begin
		isPrime = 1;
	end	else if (num==16'd42589) begin
		isPrime = 1;
	end	else if (num==16'd42611) begin
		isPrime = 1;
	end	else if (num==16'd42641) begin
		isPrime = 1;
	end	else if (num==16'd42643) begin
		isPrime = 1;
	end	else if (num==16'd42649) begin
		isPrime = 1;
	end	else if (num==16'd42667) begin
		isPrime = 1;
	end	else if (num==16'd42677) begin
		isPrime = 1;
	end	else if (num==16'd42683) begin
		isPrime = 1;
	end	else if (num==16'd42689) begin
		isPrime = 1;
	end	else if (num==16'd42697) begin
		isPrime = 1;
	end	else if (num==16'd42701) begin
		isPrime = 1;
	end	else if (num==16'd42703) begin
		isPrime = 1;
	end	else if (num==16'd42709) begin
		isPrime = 1;
	end	else if (num==16'd42719) begin
		isPrime = 1;
	end	else if (num==16'd42727) begin
		isPrime = 1;
	end	else if (num==16'd42737) begin
		isPrime = 1;
	end	else if (num==16'd42743) begin
		isPrime = 1;
	end	else if (num==16'd42751) begin
		isPrime = 1;
	end	else if (num==16'd42767) begin
		isPrime = 1;
	end	else if (num==16'd42773) begin
		isPrime = 1;
	end	else if (num==16'd42787) begin
		isPrime = 1;
	end	else if (num==16'd42793) begin
		isPrime = 1;
	end	else if (num==16'd42797) begin
		isPrime = 1;
	end	else if (num==16'd42821) begin
		isPrime = 1;
	end	else if (num==16'd42829) begin
		isPrime = 1;
	end	else if (num==16'd42839) begin
		isPrime = 1;
	end	else if (num==16'd42841) begin
		isPrime = 1;
	end	else if (num==16'd42853) begin
		isPrime = 1;
	end	else if (num==16'd42859) begin
		isPrime = 1;
	end	else if (num==16'd42863) begin
		isPrime = 1;
	end	else if (num==16'd42899) begin
		isPrime = 1;
	end	else if (num==16'd42901) begin
		isPrime = 1;
	end	else if (num==16'd42923) begin
		isPrime = 1;
	end	else if (num==16'd42929) begin
		isPrime = 1;
	end	else if (num==16'd42937) begin
		isPrime = 1;
	end	else if (num==16'd42943) begin
		isPrime = 1;
	end	else if (num==16'd42953) begin
		isPrime = 1;
	end	else if (num==16'd42961) begin
		isPrime = 1;
	end	else if (num==16'd42967) begin
		isPrime = 1;
	end	else if (num==16'd42979) begin
		isPrime = 1;
	end	else if (num==16'd42989) begin
		isPrime = 1;
	end	else if (num==16'd43003) begin
		isPrime = 1;
	end	else if (num==16'd43013) begin
		isPrime = 1;
	end	else if (num==16'd43019) begin
		isPrime = 1;
	end	else if (num==16'd43037) begin
		isPrime = 1;
	end	else if (num==16'd43049) begin
		isPrime = 1;
	end	else if (num==16'd43051) begin
		isPrime = 1;
	end	else if (num==16'd43063) begin
		isPrime = 1;
	end	else if (num==16'd43067) begin
		isPrime = 1;
	end	else if (num==16'd43093) begin
		isPrime = 1;
	end	else if (num==16'd43103) begin
		isPrime = 1;
	end	else if (num==16'd43117) begin
		isPrime = 1;
	end	else if (num==16'd43133) begin
		isPrime = 1;
	end	else if (num==16'd43151) begin
		isPrime = 1;
	end	else if (num==16'd43159) begin
		isPrime = 1;
	end	else if (num==16'd43177) begin
		isPrime = 1;
	end	else if (num==16'd43189) begin
		isPrime = 1;
	end	else if (num==16'd43201) begin
		isPrime = 1;
	end	else if (num==16'd43207) begin
		isPrime = 1;
	end	else if (num==16'd43223) begin
		isPrime = 1;
	end	else if (num==16'd43237) begin
		isPrime = 1;
	end	else if (num==16'd43261) begin
		isPrime = 1;
	end	else if (num==16'd43271) begin
		isPrime = 1;
	end	else if (num==16'd43283) begin
		isPrime = 1;
	end	else if (num==16'd43291) begin
		isPrime = 1;
	end	else if (num==16'd43313) begin
		isPrime = 1;
	end	else if (num==16'd43319) begin
		isPrime = 1;
	end	else if (num==16'd43321) begin
		isPrime = 1;
	end	else if (num==16'd43331) begin
		isPrime = 1;
	end	else if (num==16'd43391) begin
		isPrime = 1;
	end	else if (num==16'd43397) begin
		isPrime = 1;
	end	else if (num==16'd43399) begin
		isPrime = 1;
	end	else if (num==16'd43403) begin
		isPrime = 1;
	end	else if (num==16'd43411) begin
		isPrime = 1;
	end	else if (num==16'd43427) begin
		isPrime = 1;
	end	else if (num==16'd43441) begin
		isPrime = 1;
	end	else if (num==16'd43451) begin
		isPrime = 1;
	end	else if (num==16'd43457) begin
		isPrime = 1;
	end	else if (num==16'd43481) begin
		isPrime = 1;
	end	else if (num==16'd43487) begin
		isPrime = 1;
	end	else if (num==16'd43499) begin
		isPrime = 1;
	end	else if (num==16'd43517) begin
		isPrime = 1;
	end	else if (num==16'd43541) begin
		isPrime = 1;
	end	else if (num==16'd43543) begin
		isPrime = 1;
	end	else if (num==16'd43573) begin
		isPrime = 1;
	end	else if (num==16'd43577) begin
		isPrime = 1;
	end	else if (num==16'd43579) begin
		isPrime = 1;
	end	else if (num==16'd43591) begin
		isPrime = 1;
	end	else if (num==16'd43597) begin
		isPrime = 1;
	end	else if (num==16'd43607) begin
		isPrime = 1;
	end	else if (num==16'd43609) begin
		isPrime = 1;
	end	else if (num==16'd43613) begin
		isPrime = 1;
	end	else if (num==16'd43627) begin
		isPrime = 1;
	end	else if (num==16'd43633) begin
		isPrime = 1;
	end	else if (num==16'd43649) begin
		isPrime = 1;
	end	else if (num==16'd43651) begin
		isPrime = 1;
	end	else if (num==16'd43661) begin
		isPrime = 1;
	end	else if (num==16'd43669) begin
		isPrime = 1;
	end	else if (num==16'd43691) begin
		isPrime = 1;
	end	else if (num==16'd43711) begin
		isPrime = 1;
	end	else if (num==16'd43717) begin
		isPrime = 1;
	end	else if (num==16'd43721) begin
		isPrime = 1;
	end	else if (num==16'd43753) begin
		isPrime = 1;
	end	else if (num==16'd43759) begin
		isPrime = 1;
	end	else if (num==16'd43777) begin
		isPrime = 1;
	end	else if (num==16'd43781) begin
		isPrime = 1;
	end	else if (num==16'd43783) begin
		isPrime = 1;
	end	else if (num==16'd43787) begin
		isPrime = 1;
	end	else if (num==16'd43789) begin
		isPrime = 1;
	end	else if (num==16'd43793) begin
		isPrime = 1;
	end	else if (num==16'd43801) begin
		isPrime = 1;
	end	else if (num==16'd43853) begin
		isPrime = 1;
	end	else if (num==16'd43867) begin
		isPrime = 1;
	end	else if (num==16'd43889) begin
		isPrime = 1;
	end	else if (num==16'd43891) begin
		isPrime = 1;
	end	else if (num==16'd43913) begin
		isPrime = 1;
	end	else if (num==16'd43933) begin
		isPrime = 1;
	end	else if (num==16'd43943) begin
		isPrime = 1;
	end	else if (num==16'd43951) begin
		isPrime = 1;
	end	else if (num==16'd43961) begin
		isPrime = 1;
	end	else if (num==16'd43963) begin
		isPrime = 1;
	end	else if (num==16'd43969) begin
		isPrime = 1;
	end	else if (num==16'd43973) begin
		isPrime = 1;
	end	else if (num==16'd43987) begin
		isPrime = 1;
	end	else if (num==16'd43991) begin
		isPrime = 1;
	end	else if (num==16'd43997) begin
		isPrime = 1;
	end	else if (num==16'd44017) begin
		isPrime = 1;
	end	else if (num==16'd44021) begin
		isPrime = 1;
	end	else if (num==16'd44027) begin
		isPrime = 1;
	end	else if (num==16'd44029) begin
		isPrime = 1;
	end	else if (num==16'd44041) begin
		isPrime = 1;
	end	else if (num==16'd44053) begin
		isPrime = 1;
	end	else if (num==16'd44059) begin
		isPrime = 1;
	end	else if (num==16'd44071) begin
		isPrime = 1;
	end	else if (num==16'd44087) begin
		isPrime = 1;
	end	else if (num==16'd44089) begin
		isPrime = 1;
	end	else if (num==16'd44101) begin
		isPrime = 1;
	end	else if (num==16'd44111) begin
		isPrime = 1;
	end	else if (num==16'd44119) begin
		isPrime = 1;
	end	else if (num==16'd44123) begin
		isPrime = 1;
	end	else if (num==16'd44129) begin
		isPrime = 1;
	end	else if (num==16'd44131) begin
		isPrime = 1;
	end	else if (num==16'd44159) begin
		isPrime = 1;
	end	else if (num==16'd44171) begin
		isPrime = 1;
	end	else if (num==16'd44179) begin
		isPrime = 1;
	end	else if (num==16'd44189) begin
		isPrime = 1;
	end	else if (num==16'd44201) begin
		isPrime = 1;
	end	else if (num==16'd44203) begin
		isPrime = 1;
	end	else if (num==16'd44207) begin
		isPrime = 1;
	end	else if (num==16'd44221) begin
		isPrime = 1;
	end	else if (num==16'd44249) begin
		isPrime = 1;
	end	else if (num==16'd44257) begin
		isPrime = 1;
	end	else if (num==16'd44263) begin
		isPrime = 1;
	end	else if (num==16'd44267) begin
		isPrime = 1;
	end	else if (num==16'd44269) begin
		isPrime = 1;
	end	else if (num==16'd44273) begin
		isPrime = 1;
	end	else if (num==16'd44279) begin
		isPrime = 1;
	end	else if (num==16'd44281) begin
		isPrime = 1;
	end	else if (num==16'd44293) begin
		isPrime = 1;
	end	else if (num==16'd44351) begin
		isPrime = 1;
	end	else if (num==16'd44357) begin
		isPrime = 1;
	end	else if (num==16'd44371) begin
		isPrime = 1;
	end	else if (num==16'd44381) begin
		isPrime = 1;
	end	else if (num==16'd44383) begin
		isPrime = 1;
	end	else if (num==16'd44389) begin
		isPrime = 1;
	end	else if (num==16'd44417) begin
		isPrime = 1;
	end	else if (num==16'd44449) begin
		isPrime = 1;
	end	else if (num==16'd44453) begin
		isPrime = 1;
	end	else if (num==16'd44483) begin
		isPrime = 1;
	end	else if (num==16'd44491) begin
		isPrime = 1;
	end	else if (num==16'd44497) begin
		isPrime = 1;
	end	else if (num==16'd44501) begin
		isPrime = 1;
	end	else if (num==16'd44507) begin
		isPrime = 1;
	end	else if (num==16'd44519) begin
		isPrime = 1;
	end	else if (num==16'd44531) begin
		isPrime = 1;
	end	else if (num==16'd44533) begin
		isPrime = 1;
	end	else if (num==16'd44537) begin
		isPrime = 1;
	end	else if (num==16'd44543) begin
		isPrime = 1;
	end	else if (num==16'd44549) begin
		isPrime = 1;
	end	else if (num==16'd44563) begin
		isPrime = 1;
	end	else if (num==16'd44579) begin
		isPrime = 1;
	end	else if (num==16'd44587) begin
		isPrime = 1;
	end	else if (num==16'd44617) begin
		isPrime = 1;
	end	else if (num==16'd44621) begin
		isPrime = 1;
	end	else if (num==16'd44623) begin
		isPrime = 1;
	end	else if (num==16'd44633) begin
		isPrime = 1;
	end	else if (num==16'd44641) begin
		isPrime = 1;
	end	else if (num==16'd44647) begin
		isPrime = 1;
	end	else if (num==16'd44651) begin
		isPrime = 1;
	end	else if (num==16'd44657) begin
		isPrime = 1;
	end	else if (num==16'd44683) begin
		isPrime = 1;
	end	else if (num==16'd44687) begin
		isPrime = 1;
	end	else if (num==16'd44699) begin
		isPrime = 1;
	end	else if (num==16'd44701) begin
		isPrime = 1;
	end	else if (num==16'd44711) begin
		isPrime = 1;
	end	else if (num==16'd44729) begin
		isPrime = 1;
	end	else if (num==16'd44741) begin
		isPrime = 1;
	end	else if (num==16'd44753) begin
		isPrime = 1;
	end	else if (num==16'd44771) begin
		isPrime = 1;
	end	else if (num==16'd44773) begin
		isPrime = 1;
	end	else if (num==16'd44777) begin
		isPrime = 1;
	end	else if (num==16'd44789) begin
		isPrime = 1;
	end	else if (num==16'd44797) begin
		isPrime = 1;
	end	else if (num==16'd44809) begin
		isPrime = 1;
	end	else if (num==16'd44819) begin
		isPrime = 1;
	end	else if (num==16'd44839) begin
		isPrime = 1;
	end	else if (num==16'd44843) begin
		isPrime = 1;
	end	else if (num==16'd44851) begin
		isPrime = 1;
	end	else if (num==16'd44867) begin
		isPrime = 1;
	end	else if (num==16'd44879) begin
		isPrime = 1;
	end	else if (num==16'd44887) begin
		isPrime = 1;
	end	else if (num==16'd44893) begin
		isPrime = 1;
	end	else if (num==16'd44909) begin
		isPrime = 1;
	end	else if (num==16'd44917) begin
		isPrime = 1;
	end	else if (num==16'd44927) begin
		isPrime = 1;
	end	else if (num==16'd44939) begin
		isPrime = 1;
	end	else if (num==16'd44953) begin
		isPrime = 1;
	end	else if (num==16'd44959) begin
		isPrime = 1;
	end	else if (num==16'd44963) begin
		isPrime = 1;
	end	else if (num==16'd44971) begin
		isPrime = 1;
	end	else if (num==16'd44983) begin
		isPrime = 1;
	end	else if (num==16'd44987) begin
		isPrime = 1;
	end	else if (num==16'd45007) begin
		isPrime = 1;
	end	else if (num==16'd45013) begin
		isPrime = 1;
	end	else if (num==16'd45053) begin
		isPrime = 1;
	end	else if (num==16'd45061) begin
		isPrime = 1;
	end	else if (num==16'd45077) begin
		isPrime = 1;
	end	else if (num==16'd45083) begin
		isPrime = 1;
	end	else if (num==16'd45119) begin
		isPrime = 1;
	end	else if (num==16'd45121) begin
		isPrime = 1;
	end	else if (num==16'd45127) begin
		isPrime = 1;
	end	else if (num==16'd45131) begin
		isPrime = 1;
	end	else if (num==16'd45137) begin
		isPrime = 1;
	end	else if (num==16'd45139) begin
		isPrime = 1;
	end	else if (num==16'd45161) begin
		isPrime = 1;
	end	else if (num==16'd45179) begin
		isPrime = 1;
	end	else if (num==16'd45181) begin
		isPrime = 1;
	end	else if (num==16'd45191) begin
		isPrime = 1;
	end	else if (num==16'd45197) begin
		isPrime = 1;
	end	else if (num==16'd45233) begin
		isPrime = 1;
	end	else if (num==16'd45247) begin
		isPrime = 1;
	end	else if (num==16'd45259) begin
		isPrime = 1;
	end	else if (num==16'd45263) begin
		isPrime = 1;
	end	else if (num==16'd45281) begin
		isPrime = 1;
	end	else if (num==16'd45289) begin
		isPrime = 1;
	end	else if (num==16'd45293) begin
		isPrime = 1;
	end	else if (num==16'd45307) begin
		isPrime = 1;
	end	else if (num==16'd45317) begin
		isPrime = 1;
	end	else if (num==16'd45319) begin
		isPrime = 1;
	end	else if (num==16'd45329) begin
		isPrime = 1;
	end	else if (num==16'd45337) begin
		isPrime = 1;
	end	else if (num==16'd45341) begin
		isPrime = 1;
	end	else if (num==16'd45343) begin
		isPrime = 1;
	end	else if (num==16'd45361) begin
		isPrime = 1;
	end	else if (num==16'd45377) begin
		isPrime = 1;
	end	else if (num==16'd45389) begin
		isPrime = 1;
	end	else if (num==16'd45403) begin
		isPrime = 1;
	end	else if (num==16'd45413) begin
		isPrime = 1;
	end	else if (num==16'd45427) begin
		isPrime = 1;
	end	else if (num==16'd45433) begin
		isPrime = 1;
	end	else if (num==16'd45439) begin
		isPrime = 1;
	end	else if (num==16'd45481) begin
		isPrime = 1;
	end	else if (num==16'd45491) begin
		isPrime = 1;
	end	else if (num==16'd45497) begin
		isPrime = 1;
	end	else if (num==16'd45503) begin
		isPrime = 1;
	end	else if (num==16'd45523) begin
		isPrime = 1;
	end	else if (num==16'd45533) begin
		isPrime = 1;
	end	else if (num==16'd45541) begin
		isPrime = 1;
	end	else if (num==16'd45553) begin
		isPrime = 1;
	end	else if (num==16'd45557) begin
		isPrime = 1;
	end	else if (num==16'd45569) begin
		isPrime = 1;
	end	else if (num==16'd45587) begin
		isPrime = 1;
	end	else if (num==16'd45589) begin
		isPrime = 1;
	end	else if (num==16'd45599) begin
		isPrime = 1;
	end	else if (num==16'd45613) begin
		isPrime = 1;
	end	else if (num==16'd45631) begin
		isPrime = 1;
	end	else if (num==16'd45641) begin
		isPrime = 1;
	end	else if (num==16'd45659) begin
		isPrime = 1;
	end	else if (num==16'd45667) begin
		isPrime = 1;
	end	else if (num==16'd45673) begin
		isPrime = 1;
	end	else if (num==16'd45677) begin
		isPrime = 1;
	end	else if (num==16'd45691) begin
		isPrime = 1;
	end	else if (num==16'd45697) begin
		isPrime = 1;
	end	else if (num==16'd45707) begin
		isPrime = 1;
	end	else if (num==16'd45737) begin
		isPrime = 1;
	end	else if (num==16'd45751) begin
		isPrime = 1;
	end	else if (num==16'd45757) begin
		isPrime = 1;
	end	else if (num==16'd45763) begin
		isPrime = 1;
	end	else if (num==16'd45767) begin
		isPrime = 1;
	end	else if (num==16'd45779) begin
		isPrime = 1;
	end	else if (num==16'd45817) begin
		isPrime = 1;
	end	else if (num==16'd45821) begin
		isPrime = 1;
	end	else if (num==16'd45823) begin
		isPrime = 1;
	end	else if (num==16'd45827) begin
		isPrime = 1;
	end	else if (num==16'd45833) begin
		isPrime = 1;
	end	else if (num==16'd45841) begin
		isPrime = 1;
	end	else if (num==16'd45853) begin
		isPrime = 1;
	end	else if (num==16'd45863) begin
		isPrime = 1;
	end	else if (num==16'd45869) begin
		isPrime = 1;
	end	else if (num==16'd45887) begin
		isPrime = 1;
	end	else if (num==16'd45893) begin
		isPrime = 1;
	end	else if (num==16'd45943) begin
		isPrime = 1;
	end	else if (num==16'd45949) begin
		isPrime = 1;
	end	else if (num==16'd45953) begin
		isPrime = 1;
	end	else if (num==16'd45959) begin
		isPrime = 1;
	end	else if (num==16'd45971) begin
		isPrime = 1;
	end	else if (num==16'd45979) begin
		isPrime = 1;
	end	else if (num==16'd45989) begin
		isPrime = 1;
	end	else if (num==16'd46021) begin
		isPrime = 1;
	end	else if (num==16'd46027) begin
		isPrime = 1;
	end	else if (num==16'd46049) begin
		isPrime = 1;
	end	else if (num==16'd46051) begin
		isPrime = 1;
	end	else if (num==16'd46061) begin
		isPrime = 1;
	end	else if (num==16'd46073) begin
		isPrime = 1;
	end	else if (num==16'd46091) begin
		isPrime = 1;
	end	else if (num==16'd46093) begin
		isPrime = 1;
	end	else if (num==16'd46099) begin
		isPrime = 1;
	end	else if (num==16'd46103) begin
		isPrime = 1;
	end	else if (num==16'd46133) begin
		isPrime = 1;
	end	else if (num==16'd46141) begin
		isPrime = 1;
	end	else if (num==16'd46147) begin
		isPrime = 1;
	end	else if (num==16'd46153) begin
		isPrime = 1;
	end	else if (num==16'd46171) begin
		isPrime = 1;
	end	else if (num==16'd46181) begin
		isPrime = 1;
	end	else if (num==16'd46183) begin
		isPrime = 1;
	end	else if (num==16'd46187) begin
		isPrime = 1;
	end	else if (num==16'd46199) begin
		isPrime = 1;
	end	else if (num==16'd46219) begin
		isPrime = 1;
	end	else if (num==16'd46229) begin
		isPrime = 1;
	end	else if (num==16'd46237) begin
		isPrime = 1;
	end	else if (num==16'd46261) begin
		isPrime = 1;
	end	else if (num==16'd46271) begin
		isPrime = 1;
	end	else if (num==16'd46273) begin
		isPrime = 1;
	end	else if (num==16'd46279) begin
		isPrime = 1;
	end	else if (num==16'd46301) begin
		isPrime = 1;
	end	else if (num==16'd46307) begin
		isPrime = 1;
	end	else if (num==16'd46309) begin
		isPrime = 1;
	end	else if (num==16'd46327) begin
		isPrime = 1;
	end	else if (num==16'd46337) begin
		isPrime = 1;
	end	else if (num==16'd46349) begin
		isPrime = 1;
	end	else if (num==16'd46351) begin
		isPrime = 1;
	end	else if (num==16'd46381) begin
		isPrime = 1;
	end	else if (num==16'd46399) begin
		isPrime = 1;
	end	else if (num==16'd46411) begin
		isPrime = 1;
	end	else if (num==16'd46439) begin
		isPrime = 1;
	end	else if (num==16'd46441) begin
		isPrime = 1;
	end	else if (num==16'd46447) begin
		isPrime = 1;
	end	else if (num==16'd46451) begin
		isPrime = 1;
	end	else if (num==16'd46457) begin
		isPrime = 1;
	end	else if (num==16'd46471) begin
		isPrime = 1;
	end	else if (num==16'd46477) begin
		isPrime = 1;
	end	else if (num==16'd46489) begin
		isPrime = 1;
	end	else if (num==16'd46499) begin
		isPrime = 1;
	end	else if (num==16'd46507) begin
		isPrime = 1;
	end	else if (num==16'd46511) begin
		isPrime = 1;
	end	else if (num==16'd46523) begin
		isPrime = 1;
	end	else if (num==16'd46549) begin
		isPrime = 1;
	end	else if (num==16'd46559) begin
		isPrime = 1;
	end	else if (num==16'd46567) begin
		isPrime = 1;
	end	else if (num==16'd46573) begin
		isPrime = 1;
	end	else if (num==16'd46589) begin
		isPrime = 1;
	end	else if (num==16'd46591) begin
		isPrime = 1;
	end	else if (num==16'd46601) begin
		isPrime = 1;
	end	else if (num==16'd46619) begin
		isPrime = 1;
	end	else if (num==16'd46633) begin
		isPrime = 1;
	end	else if (num==16'd46639) begin
		isPrime = 1;
	end	else if (num==16'd46643) begin
		isPrime = 1;
	end	else if (num==16'd46649) begin
		isPrime = 1;
	end	else if (num==16'd46663) begin
		isPrime = 1;
	end	else if (num==16'd46679) begin
		isPrime = 1;
	end	else if (num==16'd46681) begin
		isPrime = 1;
	end	else if (num==16'd46687) begin
		isPrime = 1;
	end	else if (num==16'd46691) begin
		isPrime = 1;
	end	else if (num==16'd46703) begin
		isPrime = 1;
	end	else if (num==16'd46723) begin
		isPrime = 1;
	end	else if (num==16'd46727) begin
		isPrime = 1;
	end	else if (num==16'd46747) begin
		isPrime = 1;
	end	else if (num==16'd46751) begin
		isPrime = 1;
	end	else if (num==16'd46757) begin
		isPrime = 1;
	end	else if (num==16'd46769) begin
		isPrime = 1;
	end	else if (num==16'd46771) begin
		isPrime = 1;
	end	else if (num==16'd46807) begin
		isPrime = 1;
	end	else if (num==16'd46811) begin
		isPrime = 1;
	end	else if (num==16'd46817) begin
		isPrime = 1;
	end	else if (num==16'd46819) begin
		isPrime = 1;
	end	else if (num==16'd46829) begin
		isPrime = 1;
	end	else if (num==16'd46831) begin
		isPrime = 1;
	end	else if (num==16'd46853) begin
		isPrime = 1;
	end	else if (num==16'd46861) begin
		isPrime = 1;
	end	else if (num==16'd46867) begin
		isPrime = 1;
	end	else if (num==16'd46877) begin
		isPrime = 1;
	end	else if (num==16'd46889) begin
		isPrime = 1;
	end	else if (num==16'd46901) begin
		isPrime = 1;
	end	else if (num==16'd46919) begin
		isPrime = 1;
	end	else if (num==16'd46933) begin
		isPrime = 1;
	end	else if (num==16'd46957) begin
		isPrime = 1;
	end	else if (num==16'd46993) begin
		isPrime = 1;
	end	else if (num==16'd46997) begin
		isPrime = 1;
	end	else if (num==16'd47017) begin
		isPrime = 1;
	end	else if (num==16'd47041) begin
		isPrime = 1;
	end	else if (num==16'd47051) begin
		isPrime = 1;
	end	else if (num==16'd47057) begin
		isPrime = 1;
	end	else if (num==16'd47059) begin
		isPrime = 1;
	end	else if (num==16'd47087) begin
		isPrime = 1;
	end	else if (num==16'd47093) begin
		isPrime = 1;
	end	else if (num==16'd47111) begin
		isPrime = 1;
	end	else if (num==16'd47119) begin
		isPrime = 1;
	end	else if (num==16'd47123) begin
		isPrime = 1;
	end	else if (num==16'd47129) begin
		isPrime = 1;
	end	else if (num==16'd47137) begin
		isPrime = 1;
	end	else if (num==16'd47143) begin
		isPrime = 1;
	end	else if (num==16'd47147) begin
		isPrime = 1;
	end	else if (num==16'd47149) begin
		isPrime = 1;
	end	else if (num==16'd47161) begin
		isPrime = 1;
	end	else if (num==16'd47189) begin
		isPrime = 1;
	end	else if (num==16'd47207) begin
		isPrime = 1;
	end	else if (num==16'd47221) begin
		isPrime = 1;
	end	else if (num==16'd47237) begin
		isPrime = 1;
	end	else if (num==16'd47251) begin
		isPrime = 1;
	end	else if (num==16'd47269) begin
		isPrime = 1;
	end	else if (num==16'd47279) begin
		isPrime = 1;
	end	else if (num==16'd47287) begin
		isPrime = 1;
	end	else if (num==16'd47293) begin
		isPrime = 1;
	end	else if (num==16'd47297) begin
		isPrime = 1;
	end	else if (num==16'd47303) begin
		isPrime = 1;
	end	else if (num==16'd47309) begin
		isPrime = 1;
	end	else if (num==16'd47317) begin
		isPrime = 1;
	end	else if (num==16'd47339) begin
		isPrime = 1;
	end	else if (num==16'd47351) begin
		isPrime = 1;
	end	else if (num==16'd47353) begin
		isPrime = 1;
	end	else if (num==16'd47363) begin
		isPrime = 1;
	end	else if (num==16'd47381) begin
		isPrime = 1;
	end	else if (num==16'd47387) begin
		isPrime = 1;
	end	else if (num==16'd47389) begin
		isPrime = 1;
	end	else if (num==16'd47407) begin
		isPrime = 1;
	end	else if (num==16'd47417) begin
		isPrime = 1;
	end	else if (num==16'd47419) begin
		isPrime = 1;
	end	else if (num==16'd47431) begin
		isPrime = 1;
	end	else if (num==16'd47441) begin
		isPrime = 1;
	end	else if (num==16'd47459) begin
		isPrime = 1;
	end	else if (num==16'd47491) begin
		isPrime = 1;
	end	else if (num==16'd47497) begin
		isPrime = 1;
	end	else if (num==16'd47501) begin
		isPrime = 1;
	end	else if (num==16'd47507) begin
		isPrime = 1;
	end	else if (num==16'd47513) begin
		isPrime = 1;
	end	else if (num==16'd47521) begin
		isPrime = 1;
	end	else if (num==16'd47527) begin
		isPrime = 1;
	end	else if (num==16'd47533) begin
		isPrime = 1;
	end	else if (num==16'd47543) begin
		isPrime = 1;
	end	else if (num==16'd47563) begin
		isPrime = 1;
	end	else if (num==16'd47569) begin
		isPrime = 1;
	end	else if (num==16'd47581) begin
		isPrime = 1;
	end	else if (num==16'd47591) begin
		isPrime = 1;
	end	else if (num==16'd47599) begin
		isPrime = 1;
	end	else if (num==16'd47609) begin
		isPrime = 1;
	end	else if (num==16'd47623) begin
		isPrime = 1;
	end	else if (num==16'd47629) begin
		isPrime = 1;
	end	else if (num==16'd47639) begin
		isPrime = 1;
	end	else if (num==16'd47653) begin
		isPrime = 1;
	end	else if (num==16'd47657) begin
		isPrime = 1;
	end	else if (num==16'd47659) begin
		isPrime = 1;
	end	else if (num==16'd47681) begin
		isPrime = 1;
	end	else if (num==16'd47699) begin
		isPrime = 1;
	end	else if (num==16'd47701) begin
		isPrime = 1;
	end	else if (num==16'd47711) begin
		isPrime = 1;
	end	else if (num==16'd47713) begin
		isPrime = 1;
	end	else if (num==16'd47717) begin
		isPrime = 1;
	end	else if (num==16'd47737) begin
		isPrime = 1;
	end	else if (num==16'd47741) begin
		isPrime = 1;
	end	else if (num==16'd47743) begin
		isPrime = 1;
	end	else if (num==16'd47777) begin
		isPrime = 1;
	end	else if (num==16'd47779) begin
		isPrime = 1;
	end	else if (num==16'd47791) begin
		isPrime = 1;
	end	else if (num==16'd47797) begin
		isPrime = 1;
	end	else if (num==16'd47807) begin
		isPrime = 1;
	end	else if (num==16'd47809) begin
		isPrime = 1;
	end	else if (num==16'd47819) begin
		isPrime = 1;
	end	else if (num==16'd47837) begin
		isPrime = 1;
	end	else if (num==16'd47843) begin
		isPrime = 1;
	end	else if (num==16'd47857) begin
		isPrime = 1;
	end	else if (num==16'd47869) begin
		isPrime = 1;
	end	else if (num==16'd47881) begin
		isPrime = 1;
	end	else if (num==16'd47903) begin
		isPrime = 1;
	end	else if (num==16'd47911) begin
		isPrime = 1;
	end	else if (num==16'd47917) begin
		isPrime = 1;
	end	else if (num==16'd47933) begin
		isPrime = 1;
	end	else if (num==16'd47939) begin
		isPrime = 1;
	end	else if (num==16'd47947) begin
		isPrime = 1;
	end	else if (num==16'd47951) begin
		isPrime = 1;
	end	else if (num==16'd47963) begin
		isPrime = 1;
	end	else if (num==16'd47969) begin
		isPrime = 1;
	end	else if (num==16'd47977) begin
		isPrime = 1;
	end	else if (num==16'd47981) begin
		isPrime = 1;
	end	else if (num==16'd48017) begin
		isPrime = 1;
	end	else if (num==16'd48023) begin
		isPrime = 1;
	end	else if (num==16'd48029) begin
		isPrime = 1;
	end	else if (num==16'd48049) begin
		isPrime = 1;
	end	else if (num==16'd48073) begin
		isPrime = 1;
	end	else if (num==16'd48079) begin
		isPrime = 1;
	end	else if (num==16'd48091) begin
		isPrime = 1;
	end	else if (num==16'd48109) begin
		isPrime = 1;
	end	else if (num==16'd48119) begin
		isPrime = 1;
	end	else if (num==16'd48121) begin
		isPrime = 1;
	end	else if (num==16'd48131) begin
		isPrime = 1;
	end	else if (num==16'd48157) begin
		isPrime = 1;
	end	else if (num==16'd48163) begin
		isPrime = 1;
	end	else if (num==16'd48179) begin
		isPrime = 1;
	end	else if (num==16'd48187) begin
		isPrime = 1;
	end	else if (num==16'd48193) begin
		isPrime = 1;
	end	else if (num==16'd48197) begin
		isPrime = 1;
	end	else if (num==16'd48221) begin
		isPrime = 1;
	end	else if (num==16'd48239) begin
		isPrime = 1;
	end	else if (num==16'd48247) begin
		isPrime = 1;
	end	else if (num==16'd48259) begin
		isPrime = 1;
	end	else if (num==16'd48271) begin
		isPrime = 1;
	end	else if (num==16'd48281) begin
		isPrime = 1;
	end	else if (num==16'd48299) begin
		isPrime = 1;
	end	else if (num==16'd48311) begin
		isPrime = 1;
	end	else if (num==16'd48313) begin
		isPrime = 1;
	end	else if (num==16'd48337) begin
		isPrime = 1;
	end	else if (num==16'd48341) begin
		isPrime = 1;
	end	else if (num==16'd48353) begin
		isPrime = 1;
	end	else if (num==16'd48371) begin
		isPrime = 1;
	end	else if (num==16'd48383) begin
		isPrime = 1;
	end	else if (num==16'd48397) begin
		isPrime = 1;
	end	else if (num==16'd48407) begin
		isPrime = 1;
	end	else if (num==16'd48409) begin
		isPrime = 1;
	end	else if (num==16'd48413) begin
		isPrime = 1;
	end	else if (num==16'd48437) begin
		isPrime = 1;
	end	else if (num==16'd48449) begin
		isPrime = 1;
	end	else if (num==16'd48463) begin
		isPrime = 1;
	end	else if (num==16'd48473) begin
		isPrime = 1;
	end	else if (num==16'd48479) begin
		isPrime = 1;
	end	else if (num==16'd48481) begin
		isPrime = 1;
	end	else if (num==16'd48487) begin
		isPrime = 1;
	end	else if (num==16'd48491) begin
		isPrime = 1;
	end	else if (num==16'd48497) begin
		isPrime = 1;
	end	else if (num==16'd48523) begin
		isPrime = 1;
	end	else if (num==16'd48527) begin
		isPrime = 1;
	end	else if (num==16'd48533) begin
		isPrime = 1;
	end	else if (num==16'd48539) begin
		isPrime = 1;
	end	else if (num==16'd48541) begin
		isPrime = 1;
	end	else if (num==16'd48563) begin
		isPrime = 1;
	end	else if (num==16'd48571) begin
		isPrime = 1;
	end	else if (num==16'd48589) begin
		isPrime = 1;
	end	else if (num==16'd48593) begin
		isPrime = 1;
	end	else if (num==16'd48611) begin
		isPrime = 1;
	end	else if (num==16'd48619) begin
		isPrime = 1;
	end	else if (num==16'd48623) begin
		isPrime = 1;
	end	else if (num==16'd48647) begin
		isPrime = 1;
	end	else if (num==16'd48649) begin
		isPrime = 1;
	end	else if (num==16'd48661) begin
		isPrime = 1;
	end	else if (num==16'd48673) begin
		isPrime = 1;
	end	else if (num==16'd48677) begin
		isPrime = 1;
	end	else if (num==16'd48679) begin
		isPrime = 1;
	end	else if (num==16'd48731) begin
		isPrime = 1;
	end	else if (num==16'd48733) begin
		isPrime = 1;
	end	else if (num==16'd48751) begin
		isPrime = 1;
	end	else if (num==16'd48757) begin
		isPrime = 1;
	end	else if (num==16'd48761) begin
		isPrime = 1;
	end	else if (num==16'd48767) begin
		isPrime = 1;
	end	else if (num==16'd48779) begin
		isPrime = 1;
	end	else if (num==16'd48781) begin
		isPrime = 1;
	end	else if (num==16'd48787) begin
		isPrime = 1;
	end	else if (num==16'd48799) begin
		isPrime = 1;
	end	else if (num==16'd48809) begin
		isPrime = 1;
	end	else if (num==16'd48817) begin
		isPrime = 1;
	end	else if (num==16'd48821) begin
		isPrime = 1;
	end	else if (num==16'd48823) begin
		isPrime = 1;
	end	else if (num==16'd48847) begin
		isPrime = 1;
	end	else if (num==16'd48857) begin
		isPrime = 1;
	end	else if (num==16'd48859) begin
		isPrime = 1;
	end	else if (num==16'd48869) begin
		isPrime = 1;
	end	else if (num==16'd48871) begin
		isPrime = 1;
	end	else if (num==16'd48883) begin
		isPrime = 1;
	end	else if (num==16'd48889) begin
		isPrime = 1;
	end	else if (num==16'd48907) begin
		isPrime = 1;
	end	else if (num==16'd48947) begin
		isPrime = 1;
	end	else if (num==16'd48953) begin
		isPrime = 1;
	end	else if (num==16'd48973) begin
		isPrime = 1;
	end	else if (num==16'd48989) begin
		isPrime = 1;
	end	else if (num==16'd48991) begin
		isPrime = 1;
	end	else if (num==16'd49003) begin
		isPrime = 1;
	end	else if (num==16'd49009) begin
		isPrime = 1;
	end	else if (num==16'd49019) begin
		isPrime = 1;
	end	else if (num==16'd49031) begin
		isPrime = 1;
	end	else if (num==16'd49033) begin
		isPrime = 1;
	end	else if (num==16'd49037) begin
		isPrime = 1;
	end	else if (num==16'd49043) begin
		isPrime = 1;
	end	else if (num==16'd49057) begin
		isPrime = 1;
	end	else if (num==16'd49069) begin
		isPrime = 1;
	end	else if (num==16'd49081) begin
		isPrime = 1;
	end	else if (num==16'd49103) begin
		isPrime = 1;
	end	else if (num==16'd49109) begin
		isPrime = 1;
	end	else if (num==16'd49117) begin
		isPrime = 1;
	end	else if (num==16'd49121) begin
		isPrime = 1;
	end	else if (num==16'd49123) begin
		isPrime = 1;
	end	else if (num==16'd49139) begin
		isPrime = 1;
	end	else if (num==16'd49157) begin
		isPrime = 1;
	end	else if (num==16'd49169) begin
		isPrime = 1;
	end	else if (num==16'd49171) begin
		isPrime = 1;
	end	else if (num==16'd49177) begin
		isPrime = 1;
	end	else if (num==16'd49193) begin
		isPrime = 1;
	end	else if (num==16'd49199) begin
		isPrime = 1;
	end	else if (num==16'd49201) begin
		isPrime = 1;
	end	else if (num==16'd49207) begin
		isPrime = 1;
	end	else if (num==16'd49211) begin
		isPrime = 1;
	end	else if (num==16'd49223) begin
		isPrime = 1;
	end	else if (num==16'd49253) begin
		isPrime = 1;
	end	else if (num==16'd49261) begin
		isPrime = 1;
	end	else if (num==16'd49277) begin
		isPrime = 1;
	end	else if (num==16'd49279) begin
		isPrime = 1;
	end	else if (num==16'd49297) begin
		isPrime = 1;
	end	else if (num==16'd49307) begin
		isPrime = 1;
	end	else if (num==16'd49331) begin
		isPrime = 1;
	end	else if (num==16'd49333) begin
		isPrime = 1;
	end	else if (num==16'd49339) begin
		isPrime = 1;
	end	else if (num==16'd49363) begin
		isPrime = 1;
	end	else if (num==16'd49367) begin
		isPrime = 1;
	end	else if (num==16'd49369) begin
		isPrime = 1;
	end	else if (num==16'd49391) begin
		isPrime = 1;
	end	else if (num==16'd49393) begin
		isPrime = 1;
	end	else if (num==16'd49409) begin
		isPrime = 1;
	end	else if (num==16'd49411) begin
		isPrime = 1;
	end	else if (num==16'd49417) begin
		isPrime = 1;
	end	else if (num==16'd49429) begin
		isPrime = 1;
	end	else if (num==16'd49433) begin
		isPrime = 1;
	end	else if (num==16'd49451) begin
		isPrime = 1;
	end	else if (num==16'd49459) begin
		isPrime = 1;
	end	else if (num==16'd49463) begin
		isPrime = 1;
	end	else if (num==16'd49477) begin
		isPrime = 1;
	end	else if (num==16'd49481) begin
		isPrime = 1;
	end	else if (num==16'd49499) begin
		isPrime = 1;
	end	else if (num==16'd49523) begin
		isPrime = 1;
	end	else if (num==16'd49529) begin
		isPrime = 1;
	end	else if (num==16'd49531) begin
		isPrime = 1;
	end	else if (num==16'd49537) begin
		isPrime = 1;
	end	else if (num==16'd49547) begin
		isPrime = 1;
	end	else if (num==16'd49549) begin
		isPrime = 1;
	end	else if (num==16'd49559) begin
		isPrime = 1;
	end	else if (num==16'd49597) begin
		isPrime = 1;
	end	else if (num==16'd49603) begin
		isPrime = 1;
	end	else if (num==16'd49613) begin
		isPrime = 1;
	end	else if (num==16'd49627) begin
		isPrime = 1;
	end	else if (num==16'd49633) begin
		isPrime = 1;
	end	else if (num==16'd49639) begin
		isPrime = 1;
	end	else if (num==16'd49663) begin
		isPrime = 1;
	end	else if (num==16'd49667) begin
		isPrime = 1;
	end	else if (num==16'd49669) begin
		isPrime = 1;
	end	else if (num==16'd49681) begin
		isPrime = 1;
	end	else if (num==16'd49697) begin
		isPrime = 1;
	end	else if (num==16'd49711) begin
		isPrime = 1;
	end	else if (num==16'd49727) begin
		isPrime = 1;
	end	else if (num==16'd49739) begin
		isPrime = 1;
	end	else if (num==16'd49741) begin
		isPrime = 1;
	end	else if (num==16'd49747) begin
		isPrime = 1;
	end	else if (num==16'd49757) begin
		isPrime = 1;
	end	else if (num==16'd49783) begin
		isPrime = 1;
	end	else if (num==16'd49787) begin
		isPrime = 1;
	end	else if (num==16'd49789) begin
		isPrime = 1;
	end	else if (num==16'd49801) begin
		isPrime = 1;
	end	else if (num==16'd49807) begin
		isPrime = 1;
	end	else if (num==16'd49811) begin
		isPrime = 1;
	end	else if (num==16'd49823) begin
		isPrime = 1;
	end	else if (num==16'd49831) begin
		isPrime = 1;
	end	else if (num==16'd49843) begin
		isPrime = 1;
	end	else if (num==16'd49853) begin
		isPrime = 1;
	end	else if (num==16'd49871) begin
		isPrime = 1;
	end	else if (num==16'd49877) begin
		isPrime = 1;
	end	else if (num==16'd49891) begin
		isPrime = 1;
	end	else if (num==16'd49919) begin
		isPrime = 1;
	end	else if (num==16'd49921) begin
		isPrime = 1;
	end	else if (num==16'd49927) begin
		isPrime = 1;
	end	else if (num==16'd49937) begin
		isPrime = 1;
	end	else if (num==16'd49939) begin
		isPrime = 1;
	end	else if (num==16'd49943) begin
		isPrime = 1;
	end	else if (num==16'd49957) begin
		isPrime = 1;
	end	else if (num==16'd49991) begin
		isPrime = 1;
	end	else if (num==16'd49993) begin
		isPrime = 1;
	end	else if (num==16'd49999) begin
		isPrime = 1;
	end	else if (num==16'd50021) begin
		isPrime = 1;
	end	else if (num==16'd50023) begin
		isPrime = 1;
	end	else if (num==16'd50033) begin
		isPrime = 1;
	end	else if (num==16'd50047) begin
		isPrime = 1;
	end	else if (num==16'd50051) begin
		isPrime = 1;
	end	else if (num==16'd50053) begin
		isPrime = 1;
	end	else if (num==16'd50069) begin
		isPrime = 1;
	end	else if (num==16'd50077) begin
		isPrime = 1;
	end	else if (num==16'd50087) begin
		isPrime = 1;
	end	else if (num==16'd50093) begin
		isPrime = 1;
	end	else if (num==16'd50101) begin
		isPrime = 1;
	end	else if (num==16'd50111) begin
		isPrime = 1;
	end	else if (num==16'd50119) begin
		isPrime = 1;
	end	else if (num==16'd50123) begin
		isPrime = 1;
	end	else if (num==16'd50129) begin
		isPrime = 1;
	end	else if (num==16'd50131) begin
		isPrime = 1;
	end	else if (num==16'd50147) begin
		isPrime = 1;
	end	else if (num==16'd50153) begin
		isPrime = 1;
	end	else if (num==16'd50159) begin
		isPrime = 1;
	end	else if (num==16'd50177) begin
		isPrime = 1;
	end	else if (num==16'd50207) begin
		isPrime = 1;
	end	else if (num==16'd50221) begin
		isPrime = 1;
	end	else if (num==16'd50227) begin
		isPrime = 1;
	end	else if (num==16'd50231) begin
		isPrime = 1;
	end	else if (num==16'd50261) begin
		isPrime = 1;
	end	else if (num==16'd50263) begin
		isPrime = 1;
	end	else if (num==16'd50273) begin
		isPrime = 1;
	end	else if (num==16'd50287) begin
		isPrime = 1;
	end	else if (num==16'd50291) begin
		isPrime = 1;
	end	else if (num==16'd50311) begin
		isPrime = 1;
	end	else if (num==16'd50321) begin
		isPrime = 1;
	end	else if (num==16'd50329) begin
		isPrime = 1;
	end	else if (num==16'd50333) begin
		isPrime = 1;
	end	else if (num==16'd50341) begin
		isPrime = 1;
	end	else if (num==16'd50359) begin
		isPrime = 1;
	end	else if (num==16'd50363) begin
		isPrime = 1;
	end	else if (num==16'd50377) begin
		isPrime = 1;
	end	else if (num==16'd50383) begin
		isPrime = 1;
	end	else if (num==16'd50387) begin
		isPrime = 1;
	end	else if (num==16'd50411) begin
		isPrime = 1;
	end	else if (num==16'd50417) begin
		isPrime = 1;
	end	else if (num==16'd50423) begin
		isPrime = 1;
	end	else if (num==16'd50441) begin
		isPrime = 1;
	end	else if (num==16'd50459) begin
		isPrime = 1;
	end	else if (num==16'd50461) begin
		isPrime = 1;
	end	else if (num==16'd50497) begin
		isPrime = 1;
	end	else if (num==16'd50503) begin
		isPrime = 1;
	end	else if (num==16'd50513) begin
		isPrime = 1;
	end	else if (num==16'd50527) begin
		isPrime = 1;
	end	else if (num==16'd50539) begin
		isPrime = 1;
	end	else if (num==16'd50543) begin
		isPrime = 1;
	end	else if (num==16'd50549) begin
		isPrime = 1;
	end	else if (num==16'd50551) begin
		isPrime = 1;
	end	else if (num==16'd50581) begin
		isPrime = 1;
	end	else if (num==16'd50587) begin
		isPrime = 1;
	end	else if (num==16'd50591) begin
		isPrime = 1;
	end	else if (num==16'd50593) begin
		isPrime = 1;
	end	else if (num==16'd50599) begin
		isPrime = 1;
	end	else if (num==16'd50627) begin
		isPrime = 1;
	end	else if (num==16'd50647) begin
		isPrime = 1;
	end	else if (num==16'd50651) begin
		isPrime = 1;
	end	else if (num==16'd50671) begin
		isPrime = 1;
	end	else if (num==16'd50683) begin
		isPrime = 1;
	end	else if (num==16'd50707) begin
		isPrime = 1;
	end	else if (num==16'd50723) begin
		isPrime = 1;
	end	else if (num==16'd50741) begin
		isPrime = 1;
	end	else if (num==16'd50753) begin
		isPrime = 1;
	end	else if (num==16'd50767) begin
		isPrime = 1;
	end	else if (num==16'd50773) begin
		isPrime = 1;
	end	else if (num==16'd50777) begin
		isPrime = 1;
	end	else if (num==16'd50789) begin
		isPrime = 1;
	end	else if (num==16'd50821) begin
		isPrime = 1;
	end	else if (num==16'd50833) begin
		isPrime = 1;
	end	else if (num==16'd50839) begin
		isPrime = 1;
	end	else if (num==16'd50849) begin
		isPrime = 1;
	end	else if (num==16'd50857) begin
		isPrime = 1;
	end	else if (num==16'd50867) begin
		isPrime = 1;
	end	else if (num==16'd50873) begin
		isPrime = 1;
	end	else if (num==16'd50891) begin
		isPrime = 1;
	end	else if (num==16'd50893) begin
		isPrime = 1;
	end	else if (num==16'd50909) begin
		isPrime = 1;
	end	else if (num==16'd50923) begin
		isPrime = 1;
	end	else if (num==16'd50929) begin
		isPrime = 1;
	end	else if (num==16'd50951) begin
		isPrime = 1;
	end	else if (num==16'd50957) begin
		isPrime = 1;
	end	else if (num==16'd50969) begin
		isPrime = 1;
	end	else if (num==16'd50971) begin
		isPrime = 1;
	end	else if (num==16'd50989) begin
		isPrime = 1;
	end	else if (num==16'd50993) begin
		isPrime = 1;
	end	else if (num==16'd51001) begin
		isPrime = 1;
	end	else if (num==16'd51031) begin
		isPrime = 1;
	end	else if (num==16'd51043) begin
		isPrime = 1;
	end	else if (num==16'd51047) begin
		isPrime = 1;
	end	else if (num==16'd51059) begin
		isPrime = 1;
	end	else if (num==16'd51061) begin
		isPrime = 1;
	end	else if (num==16'd51071) begin
		isPrime = 1;
	end	else if (num==16'd51109) begin
		isPrime = 1;
	end	else if (num==16'd51131) begin
		isPrime = 1;
	end	else if (num==16'd51133) begin
		isPrime = 1;
	end	else if (num==16'd51137) begin
		isPrime = 1;
	end	else if (num==16'd51151) begin
		isPrime = 1;
	end	else if (num==16'd51157) begin
		isPrime = 1;
	end	else if (num==16'd51169) begin
		isPrime = 1;
	end	else if (num==16'd51193) begin
		isPrime = 1;
	end	else if (num==16'd51197) begin
		isPrime = 1;
	end	else if (num==16'd51199) begin
		isPrime = 1;
	end	else if (num==16'd51203) begin
		isPrime = 1;
	end	else if (num==16'd51217) begin
		isPrime = 1;
	end	else if (num==16'd51229) begin
		isPrime = 1;
	end	else if (num==16'd51239) begin
		isPrime = 1;
	end	else if (num==16'd51241) begin
		isPrime = 1;
	end	else if (num==16'd51257) begin
		isPrime = 1;
	end	else if (num==16'd51263) begin
		isPrime = 1;
	end	else if (num==16'd51283) begin
		isPrime = 1;
	end	else if (num==16'd51287) begin
		isPrime = 1;
	end	else if (num==16'd51307) begin
		isPrime = 1;
	end	else if (num==16'd51329) begin
		isPrime = 1;
	end	else if (num==16'd51341) begin
		isPrime = 1;
	end	else if (num==16'd51343) begin
		isPrime = 1;
	end	else if (num==16'd51347) begin
		isPrime = 1;
	end	else if (num==16'd51349) begin
		isPrime = 1;
	end	else if (num==16'd51361) begin
		isPrime = 1;
	end	else if (num==16'd51383) begin
		isPrime = 1;
	end	else if (num==16'd51407) begin
		isPrime = 1;
	end	else if (num==16'd51413) begin
		isPrime = 1;
	end	else if (num==16'd51419) begin
		isPrime = 1;
	end	else if (num==16'd51421) begin
		isPrime = 1;
	end	else if (num==16'd51427) begin
		isPrime = 1;
	end	else if (num==16'd51431) begin
		isPrime = 1;
	end	else if (num==16'd51437) begin
		isPrime = 1;
	end	else if (num==16'd51439) begin
		isPrime = 1;
	end	else if (num==16'd51449) begin
		isPrime = 1;
	end	else if (num==16'd51461) begin
		isPrime = 1;
	end	else if (num==16'd51473) begin
		isPrime = 1;
	end	else if (num==16'd51479) begin
		isPrime = 1;
	end	else if (num==16'd51481) begin
		isPrime = 1;
	end	else if (num==16'd51487) begin
		isPrime = 1;
	end	else if (num==16'd51503) begin
		isPrime = 1;
	end	else if (num==16'd51511) begin
		isPrime = 1;
	end	else if (num==16'd51517) begin
		isPrime = 1;
	end	else if (num==16'd51521) begin
		isPrime = 1;
	end	else if (num==16'd51539) begin
		isPrime = 1;
	end	else if (num==16'd51551) begin
		isPrime = 1;
	end	else if (num==16'd51563) begin
		isPrime = 1;
	end	else if (num==16'd51577) begin
		isPrime = 1;
	end	else if (num==16'd51581) begin
		isPrime = 1;
	end	else if (num==16'd51593) begin
		isPrime = 1;
	end	else if (num==16'd51599) begin
		isPrime = 1;
	end	else if (num==16'd51607) begin
		isPrime = 1;
	end	else if (num==16'd51613) begin
		isPrime = 1;
	end	else if (num==16'd51631) begin
		isPrime = 1;
	end	else if (num==16'd51637) begin
		isPrime = 1;
	end	else if (num==16'd51647) begin
		isPrime = 1;
	end	else if (num==16'd51659) begin
		isPrime = 1;
	end	else if (num==16'd51673) begin
		isPrime = 1;
	end	else if (num==16'd51679) begin
		isPrime = 1;
	end	else if (num==16'd51683) begin
		isPrime = 1;
	end	else if (num==16'd51691) begin
		isPrime = 1;
	end	else if (num==16'd51713) begin
		isPrime = 1;
	end	else if (num==16'd51719) begin
		isPrime = 1;
	end	else if (num==16'd51721) begin
		isPrime = 1;
	end	else if (num==16'd51749) begin
		isPrime = 1;
	end	else if (num==16'd51767) begin
		isPrime = 1;
	end	else if (num==16'd51769) begin
		isPrime = 1;
	end	else if (num==16'd51787) begin
		isPrime = 1;
	end	else if (num==16'd51797) begin
		isPrime = 1;
	end	else if (num==16'd51803) begin
		isPrime = 1;
	end	else if (num==16'd51817) begin
		isPrime = 1;
	end	else if (num==16'd51827) begin
		isPrime = 1;
	end	else if (num==16'd51829) begin
		isPrime = 1;
	end	else if (num==16'd51839) begin
		isPrime = 1;
	end	else if (num==16'd51853) begin
		isPrime = 1;
	end	else if (num==16'd51859) begin
		isPrime = 1;
	end	else if (num==16'd51869) begin
		isPrime = 1;
	end	else if (num==16'd51871) begin
		isPrime = 1;
	end	else if (num==16'd51893) begin
		isPrime = 1;
	end	else if (num==16'd51899) begin
		isPrime = 1;
	end	else if (num==16'd51907) begin
		isPrime = 1;
	end	else if (num==16'd51913) begin
		isPrime = 1;
	end	else if (num==16'd51929) begin
		isPrime = 1;
	end	else if (num==16'd51941) begin
		isPrime = 1;
	end	else if (num==16'd51949) begin
		isPrime = 1;
	end	else if (num==16'd51971) begin
		isPrime = 1;
	end	else if (num==16'd51973) begin
		isPrime = 1;
	end	else if (num==16'd51977) begin
		isPrime = 1;
	end	else if (num==16'd51991) begin
		isPrime = 1;
	end	else if (num==16'd52009) begin
		isPrime = 1;
	end	else if (num==16'd52021) begin
		isPrime = 1;
	end	else if (num==16'd52027) begin
		isPrime = 1;
	end	else if (num==16'd52051) begin
		isPrime = 1;
	end	else if (num==16'd52057) begin
		isPrime = 1;
	end	else if (num==16'd52067) begin
		isPrime = 1;
	end	else if (num==16'd52069) begin
		isPrime = 1;
	end	else if (num==16'd52081) begin
		isPrime = 1;
	end	else if (num==16'd52103) begin
		isPrime = 1;
	end	else if (num==16'd52121) begin
		isPrime = 1;
	end	else if (num==16'd52127) begin
		isPrime = 1;
	end	else if (num==16'd52147) begin
		isPrime = 1;
	end	else if (num==16'd52153) begin
		isPrime = 1;
	end	else if (num==16'd52163) begin
		isPrime = 1;
	end	else if (num==16'd52177) begin
		isPrime = 1;
	end	else if (num==16'd52181) begin
		isPrime = 1;
	end	else if (num==16'd52183) begin
		isPrime = 1;
	end	else if (num==16'd52189) begin
		isPrime = 1;
	end	else if (num==16'd52201) begin
		isPrime = 1;
	end	else if (num==16'd52223) begin
		isPrime = 1;
	end	else if (num==16'd52237) begin
		isPrime = 1;
	end	else if (num==16'd52249) begin
		isPrime = 1;
	end	else if (num==16'd52253) begin
		isPrime = 1;
	end	else if (num==16'd52259) begin
		isPrime = 1;
	end	else if (num==16'd52267) begin
		isPrime = 1;
	end	else if (num==16'd52289) begin
		isPrime = 1;
	end	else if (num==16'd52291) begin
		isPrime = 1;
	end	else if (num==16'd52301) begin
		isPrime = 1;
	end	else if (num==16'd52313) begin
		isPrime = 1;
	end	else if (num==16'd52321) begin
		isPrime = 1;
	end	else if (num==16'd52361) begin
		isPrime = 1;
	end	else if (num==16'd52363) begin
		isPrime = 1;
	end	else if (num==16'd52369) begin
		isPrime = 1;
	end	else if (num==16'd52379) begin
		isPrime = 1;
	end	else if (num==16'd52387) begin
		isPrime = 1;
	end	else if (num==16'd52391) begin
		isPrime = 1;
	end	else if (num==16'd52433) begin
		isPrime = 1;
	end	else if (num==16'd52453) begin
		isPrime = 1;
	end	else if (num==16'd52457) begin
		isPrime = 1;
	end	else if (num==16'd52489) begin
		isPrime = 1;
	end	else if (num==16'd52501) begin
		isPrime = 1;
	end	else if (num==16'd52511) begin
		isPrime = 1;
	end	else if (num==16'd52517) begin
		isPrime = 1;
	end	else if (num==16'd52529) begin
		isPrime = 1;
	end	else if (num==16'd52541) begin
		isPrime = 1;
	end	else if (num==16'd52543) begin
		isPrime = 1;
	end	else if (num==16'd52553) begin
		isPrime = 1;
	end	else if (num==16'd52561) begin
		isPrime = 1;
	end	else if (num==16'd52567) begin
		isPrime = 1;
	end	else if (num==16'd52571) begin
		isPrime = 1;
	end	else if (num==16'd52579) begin
		isPrime = 1;
	end	else if (num==16'd52583) begin
		isPrime = 1;
	end	else if (num==16'd52609) begin
		isPrime = 1;
	end	else if (num==16'd52627) begin
		isPrime = 1;
	end	else if (num==16'd52631) begin
		isPrime = 1;
	end	else if (num==16'd52639) begin
		isPrime = 1;
	end	else if (num==16'd52667) begin
		isPrime = 1;
	end	else if (num==16'd52673) begin
		isPrime = 1;
	end	else if (num==16'd52691) begin
		isPrime = 1;
	end	else if (num==16'd52697) begin
		isPrime = 1;
	end	else if (num==16'd52709) begin
		isPrime = 1;
	end	else if (num==16'd52711) begin
		isPrime = 1;
	end	else if (num==16'd52721) begin
		isPrime = 1;
	end	else if (num==16'd52727) begin
		isPrime = 1;
	end	else if (num==16'd52733) begin
		isPrime = 1;
	end	else if (num==16'd52747) begin
		isPrime = 1;
	end	else if (num==16'd52757) begin
		isPrime = 1;
	end	else if (num==16'd52769) begin
		isPrime = 1;
	end	else if (num==16'd52783) begin
		isPrime = 1;
	end	else if (num==16'd52807) begin
		isPrime = 1;
	end	else if (num==16'd52813) begin
		isPrime = 1;
	end	else if (num==16'd52817) begin
		isPrime = 1;
	end	else if (num==16'd52837) begin
		isPrime = 1;
	end	else if (num==16'd52859) begin
		isPrime = 1;
	end	else if (num==16'd52861) begin
		isPrime = 1;
	end	else if (num==16'd52879) begin
		isPrime = 1;
	end	else if (num==16'd52883) begin
		isPrime = 1;
	end	else if (num==16'd52889) begin
		isPrime = 1;
	end	else if (num==16'd52901) begin
		isPrime = 1;
	end	else if (num==16'd52903) begin
		isPrime = 1;
	end	else if (num==16'd52919) begin
		isPrime = 1;
	end	else if (num==16'd52937) begin
		isPrime = 1;
	end	else if (num==16'd52951) begin
		isPrime = 1;
	end	else if (num==16'd52957) begin
		isPrime = 1;
	end	else if (num==16'd52963) begin
		isPrime = 1;
	end	else if (num==16'd52967) begin
		isPrime = 1;
	end	else if (num==16'd52973) begin
		isPrime = 1;
	end	else if (num==16'd52981) begin
		isPrime = 1;
	end	else if (num==16'd52999) begin
		isPrime = 1;
	end	else if (num==16'd53003) begin
		isPrime = 1;
	end	else if (num==16'd53017) begin
		isPrime = 1;
	end	else if (num==16'd53047) begin
		isPrime = 1;
	end	else if (num==16'd53051) begin
		isPrime = 1;
	end	else if (num==16'd53069) begin
		isPrime = 1;
	end	else if (num==16'd53077) begin
		isPrime = 1;
	end	else if (num==16'd53087) begin
		isPrime = 1;
	end	else if (num==16'd53089) begin
		isPrime = 1;
	end	else if (num==16'd53093) begin
		isPrime = 1;
	end	else if (num==16'd53101) begin
		isPrime = 1;
	end	else if (num==16'd53113) begin
		isPrime = 1;
	end	else if (num==16'd53117) begin
		isPrime = 1;
	end	else if (num==16'd53129) begin
		isPrime = 1;
	end	else if (num==16'd53147) begin
		isPrime = 1;
	end	else if (num==16'd53149) begin
		isPrime = 1;
	end	else if (num==16'd53161) begin
		isPrime = 1;
	end	else if (num==16'd53171) begin
		isPrime = 1;
	end	else if (num==16'd53173) begin
		isPrime = 1;
	end	else if (num==16'd53189) begin
		isPrime = 1;
	end	else if (num==16'd53197) begin
		isPrime = 1;
	end	else if (num==16'd53201) begin
		isPrime = 1;
	end	else if (num==16'd53231) begin
		isPrime = 1;
	end	else if (num==16'd53233) begin
		isPrime = 1;
	end	else if (num==16'd53239) begin
		isPrime = 1;
	end	else if (num==16'd53267) begin
		isPrime = 1;
	end	else if (num==16'd53269) begin
		isPrime = 1;
	end	else if (num==16'd53279) begin
		isPrime = 1;
	end	else if (num==16'd53281) begin
		isPrime = 1;
	end	else if (num==16'd53299) begin
		isPrime = 1;
	end	else if (num==16'd53309) begin
		isPrime = 1;
	end	else if (num==16'd53323) begin
		isPrime = 1;
	end	else if (num==16'd53327) begin
		isPrime = 1;
	end	else if (num==16'd53353) begin
		isPrime = 1;
	end	else if (num==16'd53359) begin
		isPrime = 1;
	end	else if (num==16'd53377) begin
		isPrime = 1;
	end	else if (num==16'd53381) begin
		isPrime = 1;
	end	else if (num==16'd53401) begin
		isPrime = 1;
	end	else if (num==16'd53407) begin
		isPrime = 1;
	end	else if (num==16'd53411) begin
		isPrime = 1;
	end	else if (num==16'd53419) begin
		isPrime = 1;
	end	else if (num==16'd53437) begin
		isPrime = 1;
	end	else if (num==16'd53441) begin
		isPrime = 1;
	end	else if (num==16'd53453) begin
		isPrime = 1;
	end	else if (num==16'd53479) begin
		isPrime = 1;
	end	else if (num==16'd53503) begin
		isPrime = 1;
	end	else if (num==16'd53507) begin
		isPrime = 1;
	end	else if (num==16'd53527) begin
		isPrime = 1;
	end	else if (num==16'd53549) begin
		isPrime = 1;
	end	else if (num==16'd53551) begin
		isPrime = 1;
	end	else if (num==16'd53569) begin
		isPrime = 1;
	end	else if (num==16'd53591) begin
		isPrime = 1;
	end	else if (num==16'd53593) begin
		isPrime = 1;
	end	else if (num==16'd53597) begin
		isPrime = 1;
	end	else if (num==16'd53609) begin
		isPrime = 1;
	end	else if (num==16'd53611) begin
		isPrime = 1;
	end	else if (num==16'd53617) begin
		isPrime = 1;
	end	else if (num==16'd53623) begin
		isPrime = 1;
	end	else if (num==16'd53629) begin
		isPrime = 1;
	end	else if (num==16'd53633) begin
		isPrime = 1;
	end	else if (num==16'd53639) begin
		isPrime = 1;
	end	else if (num==16'd53653) begin
		isPrime = 1;
	end	else if (num==16'd53657) begin
		isPrime = 1;
	end	else if (num==16'd53681) begin
		isPrime = 1;
	end	else if (num==16'd53693) begin
		isPrime = 1;
	end	else if (num==16'd53699) begin
		isPrime = 1;
	end	else if (num==16'd53717) begin
		isPrime = 1;
	end	else if (num==16'd53719) begin
		isPrime = 1;
	end	else if (num==16'd53731) begin
		isPrime = 1;
	end	else if (num==16'd53759) begin
		isPrime = 1;
	end	else if (num==16'd53773) begin
		isPrime = 1;
	end	else if (num==16'd53777) begin
		isPrime = 1;
	end	else if (num==16'd53783) begin
		isPrime = 1;
	end	else if (num==16'd53791) begin
		isPrime = 1;
	end	else if (num==16'd53813) begin
		isPrime = 1;
	end	else if (num==16'd53819) begin
		isPrime = 1;
	end	else if (num==16'd53831) begin
		isPrime = 1;
	end	else if (num==16'd53849) begin
		isPrime = 1;
	end	else if (num==16'd53857) begin
		isPrime = 1;
	end	else if (num==16'd53861) begin
		isPrime = 1;
	end	else if (num==16'd53881) begin
		isPrime = 1;
	end	else if (num==16'd53887) begin
		isPrime = 1;
	end	else if (num==16'd53891) begin
		isPrime = 1;
	end	else if (num==16'd53897) begin
		isPrime = 1;
	end	else if (num==16'd53899) begin
		isPrime = 1;
	end	else if (num==16'd53917) begin
		isPrime = 1;
	end	else if (num==16'd53923) begin
		isPrime = 1;
	end	else if (num==16'd53927) begin
		isPrime = 1;
	end	else if (num==16'd53939) begin
		isPrime = 1;
	end	else if (num==16'd53951) begin
		isPrime = 1;
	end	else if (num==16'd53959) begin
		isPrime = 1;
	end	else if (num==16'd53987) begin
		isPrime = 1;
	end	else if (num==16'd53993) begin
		isPrime = 1;
	end	else if (num==16'd54001) begin
		isPrime = 1;
	end	else if (num==16'd54011) begin
		isPrime = 1;
	end	else if (num==16'd54013) begin
		isPrime = 1;
	end	else if (num==16'd54037) begin
		isPrime = 1;
	end	else if (num==16'd54049) begin
		isPrime = 1;
	end	else if (num==16'd54059) begin
		isPrime = 1;
	end	else if (num==16'd54083) begin
		isPrime = 1;
	end	else if (num==16'd54091) begin
		isPrime = 1;
	end	else if (num==16'd54101) begin
		isPrime = 1;
	end	else if (num==16'd54121) begin
		isPrime = 1;
	end	else if (num==16'd54133) begin
		isPrime = 1;
	end	else if (num==16'd54139) begin
		isPrime = 1;
	end	else if (num==16'd54151) begin
		isPrime = 1;
	end	else if (num==16'd54163) begin
		isPrime = 1;
	end	else if (num==16'd54167) begin
		isPrime = 1;
	end	else if (num==16'd54181) begin
		isPrime = 1;
	end	else if (num==16'd54193) begin
		isPrime = 1;
	end	else if (num==16'd54217) begin
		isPrime = 1;
	end	else if (num==16'd54251) begin
		isPrime = 1;
	end	else if (num==16'd54269) begin
		isPrime = 1;
	end	else if (num==16'd54277) begin
		isPrime = 1;
	end	else if (num==16'd54287) begin
		isPrime = 1;
	end	else if (num==16'd54293) begin
		isPrime = 1;
	end	else if (num==16'd54311) begin
		isPrime = 1;
	end	else if (num==16'd54319) begin
		isPrime = 1;
	end	else if (num==16'd54323) begin
		isPrime = 1;
	end	else if (num==16'd54331) begin
		isPrime = 1;
	end	else if (num==16'd54347) begin
		isPrime = 1;
	end	else if (num==16'd54361) begin
		isPrime = 1;
	end	else if (num==16'd54367) begin
		isPrime = 1;
	end	else if (num==16'd54371) begin
		isPrime = 1;
	end	else if (num==16'd54377) begin
		isPrime = 1;
	end	else if (num==16'd54401) begin
		isPrime = 1;
	end	else if (num==16'd54403) begin
		isPrime = 1;
	end	else if (num==16'd54409) begin
		isPrime = 1;
	end	else if (num==16'd54413) begin
		isPrime = 1;
	end	else if (num==16'd54419) begin
		isPrime = 1;
	end	else if (num==16'd54421) begin
		isPrime = 1;
	end	else if (num==16'd54437) begin
		isPrime = 1;
	end	else if (num==16'd54443) begin
		isPrime = 1;
	end	else if (num==16'd54449) begin
		isPrime = 1;
	end	else if (num==16'd54469) begin
		isPrime = 1;
	end	else if (num==16'd54493) begin
		isPrime = 1;
	end	else if (num==16'd54497) begin
		isPrime = 1;
	end	else if (num==16'd54499) begin
		isPrime = 1;
	end	else if (num==16'd54503) begin
		isPrime = 1;
	end	else if (num==16'd54517) begin
		isPrime = 1;
	end	else if (num==16'd54521) begin
		isPrime = 1;
	end	else if (num==16'd54539) begin
		isPrime = 1;
	end	else if (num==16'd54541) begin
		isPrime = 1;
	end	else if (num==16'd54547) begin
		isPrime = 1;
	end	else if (num==16'd54559) begin
		isPrime = 1;
	end	else if (num==16'd54563) begin
		isPrime = 1;
	end	else if (num==16'd54577) begin
		isPrime = 1;
	end	else if (num==16'd54581) begin
		isPrime = 1;
	end	else if (num==16'd54583) begin
		isPrime = 1;
	end	else if (num==16'd54601) begin
		isPrime = 1;
	end	else if (num==16'd54617) begin
		isPrime = 1;
	end	else if (num==16'd54623) begin
		isPrime = 1;
	end	else if (num==16'd54629) begin
		isPrime = 1;
	end	else if (num==16'd54631) begin
		isPrime = 1;
	end	else if (num==16'd54647) begin
		isPrime = 1;
	end	else if (num==16'd54667) begin
		isPrime = 1;
	end	else if (num==16'd54673) begin
		isPrime = 1;
	end	else if (num==16'd54679) begin
		isPrime = 1;
	end	else if (num==16'd54709) begin
		isPrime = 1;
	end	else if (num==16'd54713) begin
		isPrime = 1;
	end	else if (num==16'd54721) begin
		isPrime = 1;
	end	else if (num==16'd54727) begin
		isPrime = 1;
	end	else if (num==16'd54751) begin
		isPrime = 1;
	end	else if (num==16'd54767) begin
		isPrime = 1;
	end	else if (num==16'd54773) begin
		isPrime = 1;
	end	else if (num==16'd54779) begin
		isPrime = 1;
	end	else if (num==16'd54787) begin
		isPrime = 1;
	end	else if (num==16'd54799) begin
		isPrime = 1;
	end	else if (num==16'd54829) begin
		isPrime = 1;
	end	else if (num==16'd54833) begin
		isPrime = 1;
	end	else if (num==16'd54851) begin
		isPrime = 1;
	end	else if (num==16'd54869) begin
		isPrime = 1;
	end	else if (num==16'd54877) begin
		isPrime = 1;
	end	else if (num==16'd54881) begin
		isPrime = 1;
	end	else if (num==16'd54907) begin
		isPrime = 1;
	end	else if (num==16'd54917) begin
		isPrime = 1;
	end	else if (num==16'd54919) begin
		isPrime = 1;
	end	else if (num==16'd54941) begin
		isPrime = 1;
	end	else if (num==16'd54949) begin
		isPrime = 1;
	end	else if (num==16'd54959) begin
		isPrime = 1;
	end	else if (num==16'd54973) begin
		isPrime = 1;
	end	else if (num==16'd54979) begin
		isPrime = 1;
	end	else if (num==16'd54983) begin
		isPrime = 1;
	end	else if (num==16'd55001) begin
		isPrime = 1;
	end	else if (num==16'd55009) begin
		isPrime = 1;
	end	else if (num==16'd55021) begin
		isPrime = 1;
	end	else if (num==16'd55049) begin
		isPrime = 1;
	end	else if (num==16'd55051) begin
		isPrime = 1;
	end	else if (num==16'd55057) begin
		isPrime = 1;
	end	else if (num==16'd55061) begin
		isPrime = 1;
	end	else if (num==16'd55073) begin
		isPrime = 1;
	end	else if (num==16'd55079) begin
		isPrime = 1;
	end	else if (num==16'd55103) begin
		isPrime = 1;
	end	else if (num==16'd55109) begin
		isPrime = 1;
	end	else if (num==16'd55117) begin
		isPrime = 1;
	end	else if (num==16'd55127) begin
		isPrime = 1;
	end	else if (num==16'd55147) begin
		isPrime = 1;
	end	else if (num==16'd55163) begin
		isPrime = 1;
	end	else if (num==16'd55171) begin
		isPrime = 1;
	end	else if (num==16'd55201) begin
		isPrime = 1;
	end	else if (num==16'd55207) begin
		isPrime = 1;
	end	else if (num==16'd55213) begin
		isPrime = 1;
	end	else if (num==16'd55217) begin
		isPrime = 1;
	end	else if (num==16'd55219) begin
		isPrime = 1;
	end	else if (num==16'd55229) begin
		isPrime = 1;
	end	else if (num==16'd55243) begin
		isPrime = 1;
	end	else if (num==16'd55249) begin
		isPrime = 1;
	end	else if (num==16'd55259) begin
		isPrime = 1;
	end	else if (num==16'd55291) begin
		isPrime = 1;
	end	else if (num==16'd55313) begin
		isPrime = 1;
	end	else if (num==16'd55331) begin
		isPrime = 1;
	end	else if (num==16'd55333) begin
		isPrime = 1;
	end	else if (num==16'd55337) begin
		isPrime = 1;
	end	else if (num==16'd55339) begin
		isPrime = 1;
	end	else if (num==16'd55343) begin
		isPrime = 1;
	end	else if (num==16'd55351) begin
		isPrime = 1;
	end	else if (num==16'd55373) begin
		isPrime = 1;
	end	else if (num==16'd55381) begin
		isPrime = 1;
	end	else if (num==16'd55399) begin
		isPrime = 1;
	end	else if (num==16'd55411) begin
		isPrime = 1;
	end	else if (num==16'd55439) begin
		isPrime = 1;
	end	else if (num==16'd55441) begin
		isPrime = 1;
	end	else if (num==16'd55457) begin
		isPrime = 1;
	end	else if (num==16'd55469) begin
		isPrime = 1;
	end	else if (num==16'd55487) begin
		isPrime = 1;
	end	else if (num==16'd55501) begin
		isPrime = 1;
	end	else if (num==16'd55511) begin
		isPrime = 1;
	end	else if (num==16'd55529) begin
		isPrime = 1;
	end	else if (num==16'd55541) begin
		isPrime = 1;
	end	else if (num==16'd55547) begin
		isPrime = 1;
	end	else if (num==16'd55579) begin
		isPrime = 1;
	end	else if (num==16'd55589) begin
		isPrime = 1;
	end	else if (num==16'd55603) begin
		isPrime = 1;
	end	else if (num==16'd55609) begin
		isPrime = 1;
	end	else if (num==16'd55619) begin
		isPrime = 1;
	end	else if (num==16'd55621) begin
		isPrime = 1;
	end	else if (num==16'd55631) begin
		isPrime = 1;
	end	else if (num==16'd55633) begin
		isPrime = 1;
	end	else if (num==16'd55639) begin
		isPrime = 1;
	end	else if (num==16'd55661) begin
		isPrime = 1;
	end	else if (num==16'd55663) begin
		isPrime = 1;
	end	else if (num==16'd55667) begin
		isPrime = 1;
	end	else if (num==16'd55673) begin
		isPrime = 1;
	end	else if (num==16'd55681) begin
		isPrime = 1;
	end	else if (num==16'd55691) begin
		isPrime = 1;
	end	else if (num==16'd55697) begin
		isPrime = 1;
	end	else if (num==16'd55711) begin
		isPrime = 1;
	end	else if (num==16'd55717) begin
		isPrime = 1;
	end	else if (num==16'd55721) begin
		isPrime = 1;
	end	else if (num==16'd55733) begin
		isPrime = 1;
	end	else if (num==16'd55763) begin
		isPrime = 1;
	end	else if (num==16'd55787) begin
		isPrime = 1;
	end	else if (num==16'd55793) begin
		isPrime = 1;
	end	else if (num==16'd55799) begin
		isPrime = 1;
	end	else if (num==16'd55807) begin
		isPrime = 1;
	end	else if (num==16'd55813) begin
		isPrime = 1;
	end	else if (num==16'd55817) begin
		isPrime = 1;
	end	else if (num==16'd55819) begin
		isPrime = 1;
	end	else if (num==16'd55823) begin
		isPrime = 1;
	end	else if (num==16'd55829) begin
		isPrime = 1;
	end	else if (num==16'd55837) begin
		isPrime = 1;
	end	else if (num==16'd55843) begin
		isPrime = 1;
	end	else if (num==16'd55849) begin
		isPrime = 1;
	end	else if (num==16'd55871) begin
		isPrime = 1;
	end	else if (num==16'd55889) begin
		isPrime = 1;
	end	else if (num==16'd55897) begin
		isPrime = 1;
	end	else if (num==16'd55901) begin
		isPrime = 1;
	end	else if (num==16'd55903) begin
		isPrime = 1;
	end	else if (num==16'd55921) begin
		isPrime = 1;
	end	else if (num==16'd55927) begin
		isPrime = 1;
	end	else if (num==16'd55931) begin
		isPrime = 1;
	end	else if (num==16'd55933) begin
		isPrime = 1;
	end	else if (num==16'd55949) begin
		isPrime = 1;
	end	else if (num==16'd55967) begin
		isPrime = 1;
	end	else if (num==16'd55987) begin
		isPrime = 1;
	end	else if (num==16'd55997) begin
		isPrime = 1;
	end	else if (num==16'd56003) begin
		isPrime = 1;
	end	else if (num==16'd56009) begin
		isPrime = 1;
	end	else if (num==16'd56039) begin
		isPrime = 1;
	end	else if (num==16'd56041) begin
		isPrime = 1;
	end	else if (num==16'd56053) begin
		isPrime = 1;
	end	else if (num==16'd56081) begin
		isPrime = 1;
	end	else if (num==16'd56087) begin
		isPrime = 1;
	end	else if (num==16'd56093) begin
		isPrime = 1;
	end	else if (num==16'd56099) begin
		isPrime = 1;
	end	else if (num==16'd56101) begin
		isPrime = 1;
	end	else if (num==16'd56113) begin
		isPrime = 1;
	end	else if (num==16'd56123) begin
		isPrime = 1;
	end	else if (num==16'd56131) begin
		isPrime = 1;
	end	else if (num==16'd56149) begin
		isPrime = 1;
	end	else if (num==16'd56167) begin
		isPrime = 1;
	end	else if (num==16'd56171) begin
		isPrime = 1;
	end	else if (num==16'd56179) begin
		isPrime = 1;
	end	else if (num==16'd56197) begin
		isPrime = 1;
	end	else if (num==16'd56207) begin
		isPrime = 1;
	end	else if (num==16'd56209) begin
		isPrime = 1;
	end	else if (num==16'd56237) begin
		isPrime = 1;
	end	else if (num==16'd56239) begin
		isPrime = 1;
	end	else if (num==16'd56249) begin
		isPrime = 1;
	end	else if (num==16'd56263) begin
		isPrime = 1;
	end	else if (num==16'd56267) begin
		isPrime = 1;
	end	else if (num==16'd56269) begin
		isPrime = 1;
	end	else if (num==16'd56299) begin
		isPrime = 1;
	end	else if (num==16'd56311) begin
		isPrime = 1;
	end	else if (num==16'd56333) begin
		isPrime = 1;
	end	else if (num==16'd56359) begin
		isPrime = 1;
	end	else if (num==16'd56369) begin
		isPrime = 1;
	end	else if (num==16'd56377) begin
		isPrime = 1;
	end	else if (num==16'd56383) begin
		isPrime = 1;
	end	else if (num==16'd56393) begin
		isPrime = 1;
	end	else if (num==16'd56401) begin
		isPrime = 1;
	end	else if (num==16'd56417) begin
		isPrime = 1;
	end	else if (num==16'd56431) begin
		isPrime = 1;
	end	else if (num==16'd56437) begin
		isPrime = 1;
	end	else if (num==16'd56443) begin
		isPrime = 1;
	end	else if (num==16'd56453) begin
		isPrime = 1;
	end	else if (num==16'd56467) begin
		isPrime = 1;
	end	else if (num==16'd56473) begin
		isPrime = 1;
	end	else if (num==16'd56477) begin
		isPrime = 1;
	end	else if (num==16'd56479) begin
		isPrime = 1;
	end	else if (num==16'd56489) begin
		isPrime = 1;
	end	else if (num==16'd56501) begin
		isPrime = 1;
	end	else if (num==16'd56503) begin
		isPrime = 1;
	end	else if (num==16'd56509) begin
		isPrime = 1;
	end	else if (num==16'd56519) begin
		isPrime = 1;
	end	else if (num==16'd56527) begin
		isPrime = 1;
	end	else if (num==16'd56531) begin
		isPrime = 1;
	end	else if (num==16'd56533) begin
		isPrime = 1;
	end	else if (num==16'd56543) begin
		isPrime = 1;
	end	else if (num==16'd56569) begin
		isPrime = 1;
	end	else if (num==16'd56591) begin
		isPrime = 1;
	end	else if (num==16'd56597) begin
		isPrime = 1;
	end	else if (num==16'd56599) begin
		isPrime = 1;
	end	else if (num==16'd56611) begin
		isPrime = 1;
	end	else if (num==16'd56629) begin
		isPrime = 1;
	end	else if (num==16'd56633) begin
		isPrime = 1;
	end	else if (num==16'd56659) begin
		isPrime = 1;
	end	else if (num==16'd56663) begin
		isPrime = 1;
	end	else if (num==16'd56671) begin
		isPrime = 1;
	end	else if (num==16'd56681) begin
		isPrime = 1;
	end	else if (num==16'd56687) begin
		isPrime = 1;
	end	else if (num==16'd56701) begin
		isPrime = 1;
	end	else if (num==16'd56711) begin
		isPrime = 1;
	end	else if (num==16'd56713) begin
		isPrime = 1;
	end	else if (num==16'd56731) begin
		isPrime = 1;
	end	else if (num==16'd56737) begin
		isPrime = 1;
	end	else if (num==16'd56747) begin
		isPrime = 1;
	end	else if (num==16'd56767) begin
		isPrime = 1;
	end	else if (num==16'd56773) begin
		isPrime = 1;
	end	else if (num==16'd56779) begin
		isPrime = 1;
	end	else if (num==16'd56783) begin
		isPrime = 1;
	end	else if (num==16'd56807) begin
		isPrime = 1;
	end	else if (num==16'd56809) begin
		isPrime = 1;
	end	else if (num==16'd56813) begin
		isPrime = 1;
	end	else if (num==16'd56821) begin
		isPrime = 1;
	end	else if (num==16'd56827) begin
		isPrime = 1;
	end	else if (num==16'd56843) begin
		isPrime = 1;
	end	else if (num==16'd56857) begin
		isPrime = 1;
	end	else if (num==16'd56873) begin
		isPrime = 1;
	end	else if (num==16'd56891) begin
		isPrime = 1;
	end	else if (num==16'd56893) begin
		isPrime = 1;
	end	else if (num==16'd56897) begin
		isPrime = 1;
	end	else if (num==16'd56909) begin
		isPrime = 1;
	end	else if (num==16'd56911) begin
		isPrime = 1;
	end	else if (num==16'd56921) begin
		isPrime = 1;
	end	else if (num==16'd56923) begin
		isPrime = 1;
	end	else if (num==16'd56929) begin
		isPrime = 1;
	end	else if (num==16'd56941) begin
		isPrime = 1;
	end	else if (num==16'd56951) begin
		isPrime = 1;
	end	else if (num==16'd56957) begin
		isPrime = 1;
	end	else if (num==16'd56963) begin
		isPrime = 1;
	end	else if (num==16'd56983) begin
		isPrime = 1;
	end	else if (num==16'd56989) begin
		isPrime = 1;
	end	else if (num==16'd56993) begin
		isPrime = 1;
	end	else if (num==16'd56999) begin
		isPrime = 1;
	end	else if (num==16'd57037) begin
		isPrime = 1;
	end	else if (num==16'd57041) begin
		isPrime = 1;
	end	else if (num==16'd57047) begin
		isPrime = 1;
	end	else if (num==16'd57059) begin
		isPrime = 1;
	end	else if (num==16'd57073) begin
		isPrime = 1;
	end	else if (num==16'd57077) begin
		isPrime = 1;
	end	else if (num==16'd57089) begin
		isPrime = 1;
	end	else if (num==16'd57097) begin
		isPrime = 1;
	end	else if (num==16'd57107) begin
		isPrime = 1;
	end	else if (num==16'd57119) begin
		isPrime = 1;
	end	else if (num==16'd57131) begin
		isPrime = 1;
	end	else if (num==16'd57139) begin
		isPrime = 1;
	end	else if (num==16'd57143) begin
		isPrime = 1;
	end	else if (num==16'd57149) begin
		isPrime = 1;
	end	else if (num==16'd57163) begin
		isPrime = 1;
	end	else if (num==16'd57173) begin
		isPrime = 1;
	end	else if (num==16'd57179) begin
		isPrime = 1;
	end	else if (num==16'd57191) begin
		isPrime = 1;
	end	else if (num==16'd57193) begin
		isPrime = 1;
	end	else if (num==16'd57203) begin
		isPrime = 1;
	end	else if (num==16'd57221) begin
		isPrime = 1;
	end	else if (num==16'd57223) begin
		isPrime = 1;
	end	else if (num==16'd57241) begin
		isPrime = 1;
	end	else if (num==16'd57251) begin
		isPrime = 1;
	end	else if (num==16'd57259) begin
		isPrime = 1;
	end	else if (num==16'd57269) begin
		isPrime = 1;
	end	else if (num==16'd57271) begin
		isPrime = 1;
	end	else if (num==16'd57283) begin
		isPrime = 1;
	end	else if (num==16'd57287) begin
		isPrime = 1;
	end	else if (num==16'd57301) begin
		isPrime = 1;
	end	else if (num==16'd57329) begin
		isPrime = 1;
	end	else if (num==16'd57331) begin
		isPrime = 1;
	end	else if (num==16'd57347) begin
		isPrime = 1;
	end	else if (num==16'd57349) begin
		isPrime = 1;
	end	else if (num==16'd57367) begin
		isPrime = 1;
	end	else if (num==16'd57373) begin
		isPrime = 1;
	end	else if (num==16'd57383) begin
		isPrime = 1;
	end	else if (num==16'd57389) begin
		isPrime = 1;
	end	else if (num==16'd57397) begin
		isPrime = 1;
	end	else if (num==16'd57413) begin
		isPrime = 1;
	end	else if (num==16'd57427) begin
		isPrime = 1;
	end	else if (num==16'd57457) begin
		isPrime = 1;
	end	else if (num==16'd57467) begin
		isPrime = 1;
	end	else if (num==16'd57487) begin
		isPrime = 1;
	end	else if (num==16'd57493) begin
		isPrime = 1;
	end	else if (num==16'd57503) begin
		isPrime = 1;
	end	else if (num==16'd57527) begin
		isPrime = 1;
	end	else if (num==16'd57529) begin
		isPrime = 1;
	end	else if (num==16'd57557) begin
		isPrime = 1;
	end	else if (num==16'd57559) begin
		isPrime = 1;
	end	else if (num==16'd57571) begin
		isPrime = 1;
	end	else if (num==16'd57587) begin
		isPrime = 1;
	end	else if (num==16'd57593) begin
		isPrime = 1;
	end	else if (num==16'd57601) begin
		isPrime = 1;
	end	else if (num==16'd57637) begin
		isPrime = 1;
	end	else if (num==16'd57641) begin
		isPrime = 1;
	end	else if (num==16'd57649) begin
		isPrime = 1;
	end	else if (num==16'd57653) begin
		isPrime = 1;
	end	else if (num==16'd57667) begin
		isPrime = 1;
	end	else if (num==16'd57679) begin
		isPrime = 1;
	end	else if (num==16'd57689) begin
		isPrime = 1;
	end	else if (num==16'd57697) begin
		isPrime = 1;
	end	else if (num==16'd57709) begin
		isPrime = 1;
	end	else if (num==16'd57713) begin
		isPrime = 1;
	end	else if (num==16'd57719) begin
		isPrime = 1;
	end	else if (num==16'd57727) begin
		isPrime = 1;
	end	else if (num==16'd57731) begin
		isPrime = 1;
	end	else if (num==16'd57737) begin
		isPrime = 1;
	end	else if (num==16'd57751) begin
		isPrime = 1;
	end	else if (num==16'd57773) begin
		isPrime = 1;
	end	else if (num==16'd57781) begin
		isPrime = 1;
	end	else if (num==16'd57787) begin
		isPrime = 1;
	end	else if (num==16'd57791) begin
		isPrime = 1;
	end	else if (num==16'd57793) begin
		isPrime = 1;
	end	else if (num==16'd57803) begin
		isPrime = 1;
	end	else if (num==16'd57809) begin
		isPrime = 1;
	end	else if (num==16'd57829) begin
		isPrime = 1;
	end	else if (num==16'd57839) begin
		isPrime = 1;
	end	else if (num==16'd57847) begin
		isPrime = 1;
	end	else if (num==16'd57853) begin
		isPrime = 1;
	end	else if (num==16'd57859) begin
		isPrime = 1;
	end	else if (num==16'd57881) begin
		isPrime = 1;
	end	else if (num==16'd57899) begin
		isPrime = 1;
	end	else if (num==16'd57901) begin
		isPrime = 1;
	end	else if (num==16'd57917) begin
		isPrime = 1;
	end	else if (num==16'd57923) begin
		isPrime = 1;
	end	else if (num==16'd57943) begin
		isPrime = 1;
	end	else if (num==16'd57947) begin
		isPrime = 1;
	end	else if (num==16'd57973) begin
		isPrime = 1;
	end	else if (num==16'd57977) begin
		isPrime = 1;
	end	else if (num==16'd57991) begin
		isPrime = 1;
	end	else if (num==16'd58013) begin
		isPrime = 1;
	end	else if (num==16'd58027) begin
		isPrime = 1;
	end	else if (num==16'd58031) begin
		isPrime = 1;
	end	else if (num==16'd58043) begin
		isPrime = 1;
	end	else if (num==16'd58049) begin
		isPrime = 1;
	end	else if (num==16'd58057) begin
		isPrime = 1;
	end	else if (num==16'd58061) begin
		isPrime = 1;
	end	else if (num==16'd58067) begin
		isPrime = 1;
	end	else if (num==16'd58073) begin
		isPrime = 1;
	end	else if (num==16'd58099) begin
		isPrime = 1;
	end	else if (num==16'd58109) begin
		isPrime = 1;
	end	else if (num==16'd58111) begin
		isPrime = 1;
	end	else if (num==16'd58129) begin
		isPrime = 1;
	end	else if (num==16'd58147) begin
		isPrime = 1;
	end	else if (num==16'd58151) begin
		isPrime = 1;
	end	else if (num==16'd58153) begin
		isPrime = 1;
	end	else if (num==16'd58169) begin
		isPrime = 1;
	end	else if (num==16'd58171) begin
		isPrime = 1;
	end	else if (num==16'd58189) begin
		isPrime = 1;
	end	else if (num==16'd58193) begin
		isPrime = 1;
	end	else if (num==16'd58199) begin
		isPrime = 1;
	end	else if (num==16'd58207) begin
		isPrime = 1;
	end	else if (num==16'd58211) begin
		isPrime = 1;
	end	else if (num==16'd58217) begin
		isPrime = 1;
	end	else if (num==16'd58229) begin
		isPrime = 1;
	end	else if (num==16'd58231) begin
		isPrime = 1;
	end	else if (num==16'd58237) begin
		isPrime = 1;
	end	else if (num==16'd58243) begin
		isPrime = 1;
	end	else if (num==16'd58271) begin
		isPrime = 1;
	end	else if (num==16'd58309) begin
		isPrime = 1;
	end	else if (num==16'd58313) begin
		isPrime = 1;
	end	else if (num==16'd58321) begin
		isPrime = 1;
	end	else if (num==16'd58337) begin
		isPrime = 1;
	end	else if (num==16'd58363) begin
		isPrime = 1;
	end	else if (num==16'd58367) begin
		isPrime = 1;
	end	else if (num==16'd58369) begin
		isPrime = 1;
	end	else if (num==16'd58379) begin
		isPrime = 1;
	end	else if (num==16'd58391) begin
		isPrime = 1;
	end	else if (num==16'd58393) begin
		isPrime = 1;
	end	else if (num==16'd58403) begin
		isPrime = 1;
	end	else if (num==16'd58411) begin
		isPrime = 1;
	end	else if (num==16'd58417) begin
		isPrime = 1;
	end	else if (num==16'd58427) begin
		isPrime = 1;
	end	else if (num==16'd58439) begin
		isPrime = 1;
	end	else if (num==16'd58441) begin
		isPrime = 1;
	end	else if (num==16'd58451) begin
		isPrime = 1;
	end	else if (num==16'd58453) begin
		isPrime = 1;
	end	else if (num==16'd58477) begin
		isPrime = 1;
	end	else if (num==16'd58481) begin
		isPrime = 1;
	end	else if (num==16'd58511) begin
		isPrime = 1;
	end	else if (num==16'd58537) begin
		isPrime = 1;
	end	else if (num==16'd58543) begin
		isPrime = 1;
	end	else if (num==16'd58549) begin
		isPrime = 1;
	end	else if (num==16'd58567) begin
		isPrime = 1;
	end	else if (num==16'd58573) begin
		isPrime = 1;
	end	else if (num==16'd58579) begin
		isPrime = 1;
	end	else if (num==16'd58601) begin
		isPrime = 1;
	end	else if (num==16'd58603) begin
		isPrime = 1;
	end	else if (num==16'd58613) begin
		isPrime = 1;
	end	else if (num==16'd58631) begin
		isPrime = 1;
	end	else if (num==16'd58657) begin
		isPrime = 1;
	end	else if (num==16'd58661) begin
		isPrime = 1;
	end	else if (num==16'd58679) begin
		isPrime = 1;
	end	else if (num==16'd58687) begin
		isPrime = 1;
	end	else if (num==16'd58693) begin
		isPrime = 1;
	end	else if (num==16'd58699) begin
		isPrime = 1;
	end	else if (num==16'd58711) begin
		isPrime = 1;
	end	else if (num==16'd58727) begin
		isPrime = 1;
	end	else if (num==16'd58733) begin
		isPrime = 1;
	end	else if (num==16'd58741) begin
		isPrime = 1;
	end	else if (num==16'd58757) begin
		isPrime = 1;
	end	else if (num==16'd58763) begin
		isPrime = 1;
	end	else if (num==16'd58771) begin
		isPrime = 1;
	end	else if (num==16'd58787) begin
		isPrime = 1;
	end	else if (num==16'd58789) begin
		isPrime = 1;
	end	else if (num==16'd58831) begin
		isPrime = 1;
	end	else if (num==16'd58889) begin
		isPrime = 1;
	end	else if (num==16'd58897) begin
		isPrime = 1;
	end	else if (num==16'd58901) begin
		isPrime = 1;
	end	else if (num==16'd58907) begin
		isPrime = 1;
	end	else if (num==16'd58909) begin
		isPrime = 1;
	end	else if (num==16'd58913) begin
		isPrime = 1;
	end	else if (num==16'd58921) begin
		isPrime = 1;
	end	else if (num==16'd58937) begin
		isPrime = 1;
	end	else if (num==16'd58943) begin
		isPrime = 1;
	end	else if (num==16'd58963) begin
		isPrime = 1;
	end	else if (num==16'd58967) begin
		isPrime = 1;
	end	else if (num==16'd58979) begin
		isPrime = 1;
	end	else if (num==16'd58991) begin
		isPrime = 1;
	end	else if (num==16'd58997) begin
		isPrime = 1;
	end	else if (num==16'd59009) begin
		isPrime = 1;
	end	else if (num==16'd59011) begin
		isPrime = 1;
	end	else if (num==16'd59021) begin
		isPrime = 1;
	end	else if (num==16'd59023) begin
		isPrime = 1;
	end	else if (num==16'd59029) begin
		isPrime = 1;
	end	else if (num==16'd59051) begin
		isPrime = 1;
	end	else if (num==16'd59053) begin
		isPrime = 1;
	end	else if (num==16'd59063) begin
		isPrime = 1;
	end	else if (num==16'd59069) begin
		isPrime = 1;
	end	else if (num==16'd59077) begin
		isPrime = 1;
	end	else if (num==16'd59083) begin
		isPrime = 1;
	end	else if (num==16'd59093) begin
		isPrime = 1;
	end	else if (num==16'd59107) begin
		isPrime = 1;
	end	else if (num==16'd59113) begin
		isPrime = 1;
	end	else if (num==16'd59119) begin
		isPrime = 1;
	end	else if (num==16'd59123) begin
		isPrime = 1;
	end	else if (num==16'd59141) begin
		isPrime = 1;
	end	else if (num==16'd59149) begin
		isPrime = 1;
	end	else if (num==16'd59159) begin
		isPrime = 1;
	end	else if (num==16'd59167) begin
		isPrime = 1;
	end	else if (num==16'd59183) begin
		isPrime = 1;
	end	else if (num==16'd59197) begin
		isPrime = 1;
	end	else if (num==16'd59207) begin
		isPrime = 1;
	end	else if (num==16'd59209) begin
		isPrime = 1;
	end	else if (num==16'd59219) begin
		isPrime = 1;
	end	else if (num==16'd59221) begin
		isPrime = 1;
	end	else if (num==16'd59233) begin
		isPrime = 1;
	end	else if (num==16'd59239) begin
		isPrime = 1;
	end	else if (num==16'd59243) begin
		isPrime = 1;
	end	else if (num==16'd59263) begin
		isPrime = 1;
	end	else if (num==16'd59273) begin
		isPrime = 1;
	end	else if (num==16'd59281) begin
		isPrime = 1;
	end	else if (num==16'd59333) begin
		isPrime = 1;
	end	else if (num==16'd59341) begin
		isPrime = 1;
	end	else if (num==16'd59351) begin
		isPrime = 1;
	end	else if (num==16'd59357) begin
		isPrime = 1;
	end	else if (num==16'd59359) begin
		isPrime = 1;
	end	else if (num==16'd59369) begin
		isPrime = 1;
	end	else if (num==16'd59377) begin
		isPrime = 1;
	end	else if (num==16'd59387) begin
		isPrime = 1;
	end	else if (num==16'd59393) begin
		isPrime = 1;
	end	else if (num==16'd59399) begin
		isPrime = 1;
	end	else if (num==16'd59407) begin
		isPrime = 1;
	end	else if (num==16'd59417) begin
		isPrime = 1;
	end	else if (num==16'd59419) begin
		isPrime = 1;
	end	else if (num==16'd59441) begin
		isPrime = 1;
	end	else if (num==16'd59443) begin
		isPrime = 1;
	end	else if (num==16'd59447) begin
		isPrime = 1;
	end	else if (num==16'd59453) begin
		isPrime = 1;
	end	else if (num==16'd59467) begin
		isPrime = 1;
	end	else if (num==16'd59471) begin
		isPrime = 1;
	end	else if (num==16'd59473) begin
		isPrime = 1;
	end	else if (num==16'd59497) begin
		isPrime = 1;
	end	else if (num==16'd59509) begin
		isPrime = 1;
	end	else if (num==16'd59513) begin
		isPrime = 1;
	end	else if (num==16'd59539) begin
		isPrime = 1;
	end	else if (num==16'd59557) begin
		isPrime = 1;
	end	else if (num==16'd59561) begin
		isPrime = 1;
	end	else if (num==16'd59567) begin
		isPrime = 1;
	end	else if (num==16'd59581) begin
		isPrime = 1;
	end	else if (num==16'd59611) begin
		isPrime = 1;
	end	else if (num==16'd59617) begin
		isPrime = 1;
	end	else if (num==16'd59621) begin
		isPrime = 1;
	end	else if (num==16'd59627) begin
		isPrime = 1;
	end	else if (num==16'd59629) begin
		isPrime = 1;
	end	else if (num==16'd59651) begin
		isPrime = 1;
	end	else if (num==16'd59659) begin
		isPrime = 1;
	end	else if (num==16'd59663) begin
		isPrime = 1;
	end	else if (num==16'd59669) begin
		isPrime = 1;
	end	else if (num==16'd59671) begin
		isPrime = 1;
	end	else if (num==16'd59693) begin
		isPrime = 1;
	end	else if (num==16'd59699) begin
		isPrime = 1;
	end	else if (num==16'd59707) begin
		isPrime = 1;
	end	else if (num==16'd59723) begin
		isPrime = 1;
	end	else if (num==16'd59729) begin
		isPrime = 1;
	end	else if (num==16'd59743) begin
		isPrime = 1;
	end	else if (num==16'd59747) begin
		isPrime = 1;
	end	else if (num==16'd59753) begin
		isPrime = 1;
	end	else if (num==16'd59771) begin
		isPrime = 1;
	end	else if (num==16'd59779) begin
		isPrime = 1;
	end	else if (num==16'd59791) begin
		isPrime = 1;
	end	else if (num==16'd59797) begin
		isPrime = 1;
	end	else if (num==16'd59809) begin
		isPrime = 1;
	end	else if (num==16'd59833) begin
		isPrime = 1;
	end	else if (num==16'd59863) begin
		isPrime = 1;
	end	else if (num==16'd59879) begin
		isPrime = 1;
	end	else if (num==16'd59887) begin
		isPrime = 1;
	end	else if (num==16'd59921) begin
		isPrime = 1;
	end	else if (num==16'd59929) begin
		isPrime = 1;
	end	else if (num==16'd59951) begin
		isPrime = 1;
	end	else if (num==16'd59957) begin
		isPrime = 1;
	end	else if (num==16'd59971) begin
		isPrime = 1;
	end	else if (num==16'd59981) begin
		isPrime = 1;
	end	else if (num==16'd59999) begin
		isPrime = 1;
	end	else if (num==16'd60013) begin
		isPrime = 1;
	end	else if (num==16'd60017) begin
		isPrime = 1;
	end	else if (num==16'd60029) begin
		isPrime = 1;
	end	else if (num==16'd60037) begin
		isPrime = 1;
	end	else if (num==16'd60041) begin
		isPrime = 1;
	end	else if (num==16'd60077) begin
		isPrime = 1;
	end	else if (num==16'd60083) begin
		isPrime = 1;
	end	else if (num==16'd60089) begin
		isPrime = 1;
	end	else if (num==16'd60091) begin
		isPrime = 1;
	end	else if (num==16'd60101) begin
		isPrime = 1;
	end	else if (num==16'd60103) begin
		isPrime = 1;
	end	else if (num==16'd60107) begin
		isPrime = 1;
	end	else if (num==16'd60127) begin
		isPrime = 1;
	end	else if (num==16'd60133) begin
		isPrime = 1;
	end	else if (num==16'd60139) begin
		isPrime = 1;
	end	else if (num==16'd60149) begin
		isPrime = 1;
	end	else if (num==16'd60161) begin
		isPrime = 1;
	end	else if (num==16'd60167) begin
		isPrime = 1;
	end	else if (num==16'd60169) begin
		isPrime = 1;
	end	else if (num==16'd60209) begin
		isPrime = 1;
	end	else if (num==16'd60217) begin
		isPrime = 1;
	end	else if (num==16'd60223) begin
		isPrime = 1;
	end	else if (num==16'd60251) begin
		isPrime = 1;
	end	else if (num==16'd60257) begin
		isPrime = 1;
	end	else if (num==16'd60259) begin
		isPrime = 1;
	end	else if (num==16'd60271) begin
		isPrime = 1;
	end	else if (num==16'd60289) begin
		isPrime = 1;
	end	else if (num==16'd60293) begin
		isPrime = 1;
	end	else if (num==16'd60317) begin
		isPrime = 1;
	end	else if (num==16'd60331) begin
		isPrime = 1;
	end	else if (num==16'd60337) begin
		isPrime = 1;
	end	else if (num==16'd60343) begin
		isPrime = 1;
	end	else if (num==16'd60353) begin
		isPrime = 1;
	end	else if (num==16'd60373) begin
		isPrime = 1;
	end	else if (num==16'd60383) begin
		isPrime = 1;
	end	else if (num==16'd60397) begin
		isPrime = 1;
	end	else if (num==16'd60413) begin
		isPrime = 1;
	end	else if (num==16'd60427) begin
		isPrime = 1;
	end	else if (num==16'd60443) begin
		isPrime = 1;
	end	else if (num==16'd60449) begin
		isPrime = 1;
	end	else if (num==16'd60457) begin
		isPrime = 1;
	end	else if (num==16'd60493) begin
		isPrime = 1;
	end	else if (num==16'd60497) begin
		isPrime = 1;
	end	else if (num==16'd60509) begin
		isPrime = 1;
	end	else if (num==16'd60521) begin
		isPrime = 1;
	end	else if (num==16'd60527) begin
		isPrime = 1;
	end	else if (num==16'd60539) begin
		isPrime = 1;
	end	else if (num==16'd60589) begin
		isPrime = 1;
	end	else if (num==16'd60601) begin
		isPrime = 1;
	end	else if (num==16'd60607) begin
		isPrime = 1;
	end	else if (num==16'd60611) begin
		isPrime = 1;
	end	else if (num==16'd60617) begin
		isPrime = 1;
	end	else if (num==16'd60623) begin
		isPrime = 1;
	end	else if (num==16'd60631) begin
		isPrime = 1;
	end	else if (num==16'd60637) begin
		isPrime = 1;
	end	else if (num==16'd60647) begin
		isPrime = 1;
	end	else if (num==16'd60649) begin
		isPrime = 1;
	end	else if (num==16'd60659) begin
		isPrime = 1;
	end	else if (num==16'd60661) begin
		isPrime = 1;
	end	else if (num==16'd60679) begin
		isPrime = 1;
	end	else if (num==16'd60689) begin
		isPrime = 1;
	end	else if (num==16'd60703) begin
		isPrime = 1;
	end	else if (num==16'd60719) begin
		isPrime = 1;
	end	else if (num==16'd60727) begin
		isPrime = 1;
	end	else if (num==16'd60733) begin
		isPrime = 1;
	end	else if (num==16'd60737) begin
		isPrime = 1;
	end	else if (num==16'd60757) begin
		isPrime = 1;
	end	else if (num==16'd60761) begin
		isPrime = 1;
	end	else if (num==16'd60763) begin
		isPrime = 1;
	end	else if (num==16'd60773) begin
		isPrime = 1;
	end	else if (num==16'd60779) begin
		isPrime = 1;
	end	else if (num==16'd60793) begin
		isPrime = 1;
	end	else if (num==16'd60811) begin
		isPrime = 1;
	end	else if (num==16'd60821) begin
		isPrime = 1;
	end	else if (num==16'd60859) begin
		isPrime = 1;
	end	else if (num==16'd60869) begin
		isPrime = 1;
	end	else if (num==16'd60887) begin
		isPrime = 1;
	end	else if (num==16'd60889) begin
		isPrime = 1;
	end	else if (num==16'd60899) begin
		isPrime = 1;
	end	else if (num==16'd60901) begin
		isPrime = 1;
	end	else if (num==16'd60913) begin
		isPrime = 1;
	end	else if (num==16'd60917) begin
		isPrime = 1;
	end	else if (num==16'd60919) begin
		isPrime = 1;
	end	else if (num==16'd60923) begin
		isPrime = 1;
	end	else if (num==16'd60937) begin
		isPrime = 1;
	end	else if (num==16'd60943) begin
		isPrime = 1;
	end	else if (num==16'd60953) begin
		isPrime = 1;
	end	else if (num==16'd60961) begin
		isPrime = 1;
	end	else if (num==16'd61001) begin
		isPrime = 1;
	end	else if (num==16'd61007) begin
		isPrime = 1;
	end	else if (num==16'd61027) begin
		isPrime = 1;
	end	else if (num==16'd61031) begin
		isPrime = 1;
	end	else if (num==16'd61043) begin
		isPrime = 1;
	end	else if (num==16'd61051) begin
		isPrime = 1;
	end	else if (num==16'd61057) begin
		isPrime = 1;
	end	else if (num==16'd61091) begin
		isPrime = 1;
	end	else if (num==16'd61099) begin
		isPrime = 1;
	end	else if (num==16'd61121) begin
		isPrime = 1;
	end	else if (num==16'd61129) begin
		isPrime = 1;
	end	else if (num==16'd61141) begin
		isPrime = 1;
	end	else if (num==16'd61151) begin
		isPrime = 1;
	end	else if (num==16'd61153) begin
		isPrime = 1;
	end	else if (num==16'd61169) begin
		isPrime = 1;
	end	else if (num==16'd61211) begin
		isPrime = 1;
	end	else if (num==16'd61223) begin
		isPrime = 1;
	end	else if (num==16'd61231) begin
		isPrime = 1;
	end	else if (num==16'd61253) begin
		isPrime = 1;
	end	else if (num==16'd61261) begin
		isPrime = 1;
	end	else if (num==16'd61283) begin
		isPrime = 1;
	end	else if (num==16'd61291) begin
		isPrime = 1;
	end	else if (num==16'd61297) begin
		isPrime = 1;
	end	else if (num==16'd61331) begin
		isPrime = 1;
	end	else if (num==16'd61333) begin
		isPrime = 1;
	end	else if (num==16'd61339) begin
		isPrime = 1;
	end	else if (num==16'd61343) begin
		isPrime = 1;
	end	else if (num==16'd61357) begin
		isPrime = 1;
	end	else if (num==16'd61363) begin
		isPrime = 1;
	end	else if (num==16'd61379) begin
		isPrime = 1;
	end	else if (num==16'd61381) begin
		isPrime = 1;
	end	else if (num==16'd61403) begin
		isPrime = 1;
	end	else if (num==16'd61409) begin
		isPrime = 1;
	end	else if (num==16'd61417) begin
		isPrime = 1;
	end	else if (num==16'd61441) begin
		isPrime = 1;
	end	else if (num==16'd61463) begin
		isPrime = 1;
	end	else if (num==16'd61469) begin
		isPrime = 1;
	end	else if (num==16'd61471) begin
		isPrime = 1;
	end	else if (num==16'd61483) begin
		isPrime = 1;
	end	else if (num==16'd61487) begin
		isPrime = 1;
	end	else if (num==16'd61493) begin
		isPrime = 1;
	end	else if (num==16'd61507) begin
		isPrime = 1;
	end	else if (num==16'd61511) begin
		isPrime = 1;
	end	else if (num==16'd61519) begin
		isPrime = 1;
	end	else if (num==16'd61543) begin
		isPrime = 1;
	end	else if (num==16'd61547) begin
		isPrime = 1;
	end	else if (num==16'd61553) begin
		isPrime = 1;
	end	else if (num==16'd61559) begin
		isPrime = 1;
	end	else if (num==16'd61561) begin
		isPrime = 1;
	end	else if (num==16'd61583) begin
		isPrime = 1;
	end	else if (num==16'd61603) begin
		isPrime = 1;
	end	else if (num==16'd61609) begin
		isPrime = 1;
	end	else if (num==16'd61613) begin
		isPrime = 1;
	end	else if (num==16'd61627) begin
		isPrime = 1;
	end	else if (num==16'd61631) begin
		isPrime = 1;
	end	else if (num==16'd61637) begin
		isPrime = 1;
	end	else if (num==16'd61643) begin
		isPrime = 1;
	end	else if (num==16'd61651) begin
		isPrime = 1;
	end	else if (num==16'd61657) begin
		isPrime = 1;
	end	else if (num==16'd61667) begin
		isPrime = 1;
	end	else if (num==16'd61673) begin
		isPrime = 1;
	end	else if (num==16'd61681) begin
		isPrime = 1;
	end	else if (num==16'd61687) begin
		isPrime = 1;
	end	else if (num==16'd61703) begin
		isPrime = 1;
	end	else if (num==16'd61717) begin
		isPrime = 1;
	end	else if (num==16'd61723) begin
		isPrime = 1;
	end	else if (num==16'd61729) begin
		isPrime = 1;
	end	else if (num==16'd61751) begin
		isPrime = 1;
	end	else if (num==16'd61757) begin
		isPrime = 1;
	end	else if (num==16'd61781) begin
		isPrime = 1;
	end	else if (num==16'd61813) begin
		isPrime = 1;
	end	else if (num==16'd61819) begin
		isPrime = 1;
	end	else if (num==16'd61837) begin
		isPrime = 1;
	end	else if (num==16'd61843) begin
		isPrime = 1;
	end	else if (num==16'd61861) begin
		isPrime = 1;
	end	else if (num==16'd61871) begin
		isPrime = 1;
	end	else if (num==16'd61879) begin
		isPrime = 1;
	end	else if (num==16'd61909) begin
		isPrime = 1;
	end	else if (num==16'd61927) begin
		isPrime = 1;
	end	else if (num==16'd61933) begin
		isPrime = 1;
	end	else if (num==16'd61949) begin
		isPrime = 1;
	end	else if (num==16'd61961) begin
		isPrime = 1;
	end	else if (num==16'd61967) begin
		isPrime = 1;
	end	else if (num==16'd61979) begin
		isPrime = 1;
	end	else if (num==16'd61981) begin
		isPrime = 1;
	end	else if (num==16'd61987) begin
		isPrime = 1;
	end	else if (num==16'd61991) begin
		isPrime = 1;
	end	else if (num==16'd62003) begin
		isPrime = 1;
	end	else if (num==16'd62011) begin
		isPrime = 1;
	end	else if (num==16'd62017) begin
		isPrime = 1;
	end	else if (num==16'd62039) begin
		isPrime = 1;
	end	else if (num==16'd62047) begin
		isPrime = 1;
	end	else if (num==16'd62053) begin
		isPrime = 1;
	end	else if (num==16'd62057) begin
		isPrime = 1;
	end	else if (num==16'd62071) begin
		isPrime = 1;
	end	else if (num==16'd62081) begin
		isPrime = 1;
	end	else if (num==16'd62099) begin
		isPrime = 1;
	end	else if (num==16'd62119) begin
		isPrime = 1;
	end	else if (num==16'd62129) begin
		isPrime = 1;
	end	else if (num==16'd62131) begin
		isPrime = 1;
	end	else if (num==16'd62137) begin
		isPrime = 1;
	end	else if (num==16'd62141) begin
		isPrime = 1;
	end	else if (num==16'd62143) begin
		isPrime = 1;
	end	else if (num==16'd62171) begin
		isPrime = 1;
	end	else if (num==16'd62189) begin
		isPrime = 1;
	end	else if (num==16'd62191) begin
		isPrime = 1;
	end	else if (num==16'd62201) begin
		isPrime = 1;
	end	else if (num==16'd62207) begin
		isPrime = 1;
	end	else if (num==16'd62213) begin
		isPrime = 1;
	end	else if (num==16'd62219) begin
		isPrime = 1;
	end	else if (num==16'd62233) begin
		isPrime = 1;
	end	else if (num==16'd62273) begin
		isPrime = 1;
	end	else if (num==16'd62297) begin
		isPrime = 1;
	end	else if (num==16'd62299) begin
		isPrime = 1;
	end	else if (num==16'd62303) begin
		isPrime = 1;
	end	else if (num==16'd62311) begin
		isPrime = 1;
	end	else if (num==16'd62323) begin
		isPrime = 1;
	end	else if (num==16'd62327) begin
		isPrime = 1;
	end	else if (num==16'd62347) begin
		isPrime = 1;
	end	else if (num==16'd62351) begin
		isPrime = 1;
	end	else if (num==16'd62383) begin
		isPrime = 1;
	end	else if (num==16'd62401) begin
		isPrime = 1;
	end	else if (num==16'd62417) begin
		isPrime = 1;
	end	else if (num==16'd62423) begin
		isPrime = 1;
	end	else if (num==16'd62459) begin
		isPrime = 1;
	end	else if (num==16'd62467) begin
		isPrime = 1;
	end	else if (num==16'd62473) begin
		isPrime = 1;
	end	else if (num==16'd62477) begin
		isPrime = 1;
	end	else if (num==16'd62483) begin
		isPrime = 1;
	end	else if (num==16'd62497) begin
		isPrime = 1;
	end	else if (num==16'd62501) begin
		isPrime = 1;
	end	else if (num==16'd62507) begin
		isPrime = 1;
	end	else if (num==16'd62533) begin
		isPrime = 1;
	end	else if (num==16'd62539) begin
		isPrime = 1;
	end	else if (num==16'd62549) begin
		isPrime = 1;
	end	else if (num==16'd62563) begin
		isPrime = 1;
	end	else if (num==16'd62581) begin
		isPrime = 1;
	end	else if (num==16'd62591) begin
		isPrime = 1;
	end	else if (num==16'd62597) begin
		isPrime = 1;
	end	else if (num==16'd62603) begin
		isPrime = 1;
	end	else if (num==16'd62617) begin
		isPrime = 1;
	end	else if (num==16'd62627) begin
		isPrime = 1;
	end	else if (num==16'd62633) begin
		isPrime = 1;
	end	else if (num==16'd62639) begin
		isPrime = 1;
	end	else if (num==16'd62653) begin
		isPrime = 1;
	end	else if (num==16'd62659) begin
		isPrime = 1;
	end	else if (num==16'd62683) begin
		isPrime = 1;
	end	else if (num==16'd62687) begin
		isPrime = 1;
	end	else if (num==16'd62701) begin
		isPrime = 1;
	end	else if (num==16'd62723) begin
		isPrime = 1;
	end	else if (num==16'd62731) begin
		isPrime = 1;
	end	else if (num==16'd62743) begin
		isPrime = 1;
	end	else if (num==16'd62753) begin
		isPrime = 1;
	end	else if (num==16'd62761) begin
		isPrime = 1;
	end	else if (num==16'd62773) begin
		isPrime = 1;
	end	else if (num==16'd62791) begin
		isPrime = 1;
	end	else if (num==16'd62801) begin
		isPrime = 1;
	end	else if (num==16'd62819) begin
		isPrime = 1;
	end	else if (num==16'd62827) begin
		isPrime = 1;
	end	else if (num==16'd62851) begin
		isPrime = 1;
	end	else if (num==16'd62861) begin
		isPrime = 1;
	end	else if (num==16'd62869) begin
		isPrime = 1;
	end	else if (num==16'd62873) begin
		isPrime = 1;
	end	else if (num==16'd62897) begin
		isPrime = 1;
	end	else if (num==16'd62903) begin
		isPrime = 1;
	end	else if (num==16'd62921) begin
		isPrime = 1;
	end	else if (num==16'd62927) begin
		isPrime = 1;
	end	else if (num==16'd62929) begin
		isPrime = 1;
	end	else if (num==16'd62939) begin
		isPrime = 1;
	end	else if (num==16'd62969) begin
		isPrime = 1;
	end	else if (num==16'd62971) begin
		isPrime = 1;
	end	else if (num==16'd62981) begin
		isPrime = 1;
	end	else if (num==16'd62983) begin
		isPrime = 1;
	end	else if (num==16'd62987) begin
		isPrime = 1;
	end	else if (num==16'd62989) begin
		isPrime = 1;
	end	else if (num==16'd63029) begin
		isPrime = 1;
	end	else if (num==16'd63031) begin
		isPrime = 1;
	end	else if (num==16'd63059) begin
		isPrime = 1;
	end	else if (num==16'd63067) begin
		isPrime = 1;
	end	else if (num==16'd63073) begin
		isPrime = 1;
	end	else if (num==16'd63079) begin
		isPrime = 1;
	end	else if (num==16'd63097) begin
		isPrime = 1;
	end	else if (num==16'd63103) begin
		isPrime = 1;
	end	else if (num==16'd63113) begin
		isPrime = 1;
	end	else if (num==16'd63127) begin
		isPrime = 1;
	end	else if (num==16'd63131) begin
		isPrime = 1;
	end	else if (num==16'd63149) begin
		isPrime = 1;
	end	else if (num==16'd63179) begin
		isPrime = 1;
	end	else if (num==16'd63197) begin
		isPrime = 1;
	end	else if (num==16'd63199) begin
		isPrime = 1;
	end	else if (num==16'd63211) begin
		isPrime = 1;
	end	else if (num==16'd63241) begin
		isPrime = 1;
	end	else if (num==16'd63247) begin
		isPrime = 1;
	end	else if (num==16'd63277) begin
		isPrime = 1;
	end	else if (num==16'd63281) begin
		isPrime = 1;
	end	else if (num==16'd63299) begin
		isPrime = 1;
	end	else if (num==16'd63311) begin
		isPrime = 1;
	end	else if (num==16'd63313) begin
		isPrime = 1;
	end	else if (num==16'd63317) begin
		isPrime = 1;
	end	else if (num==16'd63331) begin
		isPrime = 1;
	end	else if (num==16'd63337) begin
		isPrime = 1;
	end	else if (num==16'd63347) begin
		isPrime = 1;
	end	else if (num==16'd63353) begin
		isPrime = 1;
	end	else if (num==16'd63361) begin
		isPrime = 1;
	end	else if (num==16'd63367) begin
		isPrime = 1;
	end	else if (num==16'd63377) begin
		isPrime = 1;
	end	else if (num==16'd63389) begin
		isPrime = 1;
	end	else if (num==16'd63391) begin
		isPrime = 1;
	end	else if (num==16'd63397) begin
		isPrime = 1;
	end	else if (num==16'd63409) begin
		isPrime = 1;
	end	else if (num==16'd63419) begin
		isPrime = 1;
	end	else if (num==16'd63421) begin
		isPrime = 1;
	end	else if (num==16'd63439) begin
		isPrime = 1;
	end	else if (num==16'd63443) begin
		isPrime = 1;
	end	else if (num==16'd63463) begin
		isPrime = 1;
	end	else if (num==16'd63467) begin
		isPrime = 1;
	end	else if (num==16'd63473) begin
		isPrime = 1;
	end	else if (num==16'd63487) begin
		isPrime = 1;
	end	else if (num==16'd63493) begin
		isPrime = 1;
	end	else if (num==16'd63499) begin
		isPrime = 1;
	end	else if (num==16'd63521) begin
		isPrime = 1;
	end	else if (num==16'd63527) begin
		isPrime = 1;
	end	else if (num==16'd63533) begin
		isPrime = 1;
	end	else if (num==16'd63541) begin
		isPrime = 1;
	end	else if (num==16'd63559) begin
		isPrime = 1;
	end	else if (num==16'd63577) begin
		isPrime = 1;
	end	else if (num==16'd63587) begin
		isPrime = 1;
	end	else if (num==16'd63589) begin
		isPrime = 1;
	end	else if (num==16'd63599) begin
		isPrime = 1;
	end	else if (num==16'd63601) begin
		isPrime = 1;
	end	else if (num==16'd63607) begin
		isPrime = 1;
	end	else if (num==16'd63611) begin
		isPrime = 1;
	end	else if (num==16'd63617) begin
		isPrime = 1;
	end	else if (num==16'd63629) begin
		isPrime = 1;
	end	else if (num==16'd63647) begin
		isPrime = 1;
	end	else if (num==16'd63649) begin
		isPrime = 1;
	end	else if (num==16'd63659) begin
		isPrime = 1;
	end	else if (num==16'd63667) begin
		isPrime = 1;
	end	else if (num==16'd63671) begin
		isPrime = 1;
	end	else if (num==16'd63689) begin
		isPrime = 1;
	end	else if (num==16'd63691) begin
		isPrime = 1;
	end	else if (num==16'd63697) begin
		isPrime = 1;
	end	else if (num==16'd63703) begin
		isPrime = 1;
	end	else if (num==16'd63709) begin
		isPrime = 1;
	end	else if (num==16'd63719) begin
		isPrime = 1;
	end	else if (num==16'd63727) begin
		isPrime = 1;
	end	else if (num==16'd63737) begin
		isPrime = 1;
	end	else if (num==16'd63743) begin
		isPrime = 1;
	end	else if (num==16'd63761) begin
		isPrime = 1;
	end	else if (num==16'd63773) begin
		isPrime = 1;
	end	else if (num==16'd63781) begin
		isPrime = 1;
	end	else if (num==16'd63793) begin
		isPrime = 1;
	end	else if (num==16'd63799) begin
		isPrime = 1;
	end	else if (num==16'd63803) begin
		isPrime = 1;
	end	else if (num==16'd63809) begin
		isPrime = 1;
	end	else if (num==16'd63823) begin
		isPrime = 1;
	end	else if (num==16'd63839) begin
		isPrime = 1;
	end	else if (num==16'd63841) begin
		isPrime = 1;
	end	else if (num==16'd63853) begin
		isPrime = 1;
	end	else if (num==16'd63857) begin
		isPrime = 1;
	end	else if (num==16'd63863) begin
		isPrime = 1;
	end	else if (num==16'd63901) begin
		isPrime = 1;
	end	else if (num==16'd63907) begin
		isPrime = 1;
	end	else if (num==16'd63913) begin
		isPrime = 1;
	end	else if (num==16'd63929) begin
		isPrime = 1;
	end	else if (num==16'd63949) begin
		isPrime = 1;
	end	else if (num==16'd63977) begin
		isPrime = 1;
	end	else if (num==16'd63997) begin
		isPrime = 1;
	end	else if (num==16'd64007) begin
		isPrime = 1;
	end	else if (num==16'd64013) begin
		isPrime = 1;
	end	else if (num==16'd64019) begin
		isPrime = 1;
	end	else if (num==16'd64033) begin
		isPrime = 1;
	end	else if (num==16'd64037) begin
		isPrime = 1;
	end	else if (num==16'd64063) begin
		isPrime = 1;
	end	else if (num==16'd64067) begin
		isPrime = 1;
	end	else if (num==16'd64081) begin
		isPrime = 1;
	end	else if (num==16'd64091) begin
		isPrime = 1;
	end	else if (num==16'd64109) begin
		isPrime = 1;
	end	else if (num==16'd64123) begin
		isPrime = 1;
	end	else if (num==16'd64151) begin
		isPrime = 1;
	end	else if (num==16'd64153) begin
		isPrime = 1;
	end	else if (num==16'd64157) begin
		isPrime = 1;
	end	else if (num==16'd64171) begin
		isPrime = 1;
	end	else if (num==16'd64187) begin
		isPrime = 1;
	end	else if (num==16'd64189) begin
		isPrime = 1;
	end	else if (num==16'd64217) begin
		isPrime = 1;
	end	else if (num==16'd64223) begin
		isPrime = 1;
	end	else if (num==16'd64231) begin
		isPrime = 1;
	end	else if (num==16'd64237) begin
		isPrime = 1;
	end	else if (num==16'd64271) begin
		isPrime = 1;
	end	else if (num==16'd64279) begin
		isPrime = 1;
	end	else if (num==16'd64283) begin
		isPrime = 1;
	end	else if (num==16'd64301) begin
		isPrime = 1;
	end	else if (num==16'd64303) begin
		isPrime = 1;
	end	else if (num==16'd64319) begin
		isPrime = 1;
	end	else if (num==16'd64327) begin
		isPrime = 1;
	end	else if (num==16'd64333) begin
		isPrime = 1;
	end	else if (num==16'd64373) begin
		isPrime = 1;
	end	else if (num==16'd64381) begin
		isPrime = 1;
	end	else if (num==16'd64399) begin
		isPrime = 1;
	end	else if (num==16'd64403) begin
		isPrime = 1;
	end	else if (num==16'd64433) begin
		isPrime = 1;
	end	else if (num==16'd64439) begin
		isPrime = 1;
	end	else if (num==16'd64451) begin
		isPrime = 1;
	end	else if (num==16'd64453) begin
		isPrime = 1;
	end	else if (num==16'd64483) begin
		isPrime = 1;
	end	else if (num==16'd64489) begin
		isPrime = 1;
	end	else if (num==16'd64499) begin
		isPrime = 1;
	end	else if (num==16'd64513) begin
		isPrime = 1;
	end	else if (num==16'd64553) begin
		isPrime = 1;
	end	else if (num==16'd64567) begin
		isPrime = 1;
	end	else if (num==16'd64577) begin
		isPrime = 1;
	end	else if (num==16'd64579) begin
		isPrime = 1;
	end	else if (num==16'd64591) begin
		isPrime = 1;
	end	else if (num==16'd64601) begin
		isPrime = 1;
	end	else if (num==16'd64609) begin
		isPrime = 1;
	end	else if (num==16'd64613) begin
		isPrime = 1;
	end	else if (num==16'd64621) begin
		isPrime = 1;
	end	else if (num==16'd64627) begin
		isPrime = 1;
	end	else if (num==16'd64633) begin
		isPrime = 1;
	end	else if (num==16'd64661) begin
		isPrime = 1;
	end	else if (num==16'd64663) begin
		isPrime = 1;
	end	else if (num==16'd64667) begin
		isPrime = 1;
	end	else if (num==16'd64679) begin
		isPrime = 1;
	end	else if (num==16'd64693) begin
		isPrime = 1;
	end	else if (num==16'd64709) begin
		isPrime = 1;
	end	else if (num==16'd64717) begin
		isPrime = 1;
	end	else if (num==16'd64747) begin
		isPrime = 1;
	end	else if (num==16'd64763) begin
		isPrime = 1;
	end	else if (num==16'd64781) begin
		isPrime = 1;
	end	else if (num==16'd64783) begin
		isPrime = 1;
	end	else if (num==16'd64793) begin
		isPrime = 1;
	end	else if (num==16'd64811) begin
		isPrime = 1;
	end	else if (num==16'd64817) begin
		isPrime = 1;
	end	else if (num==16'd64849) begin
		isPrime = 1;
	end	else if (num==16'd64853) begin
		isPrime = 1;
	end	else if (num==16'd64871) begin
		isPrime = 1;
	end	else if (num==16'd64877) begin
		isPrime = 1;
	end	else if (num==16'd64879) begin
		isPrime = 1;
	end	else if (num==16'd64891) begin
		isPrime = 1;
	end	else if (num==16'd64901) begin
		isPrime = 1;
	end	else if (num==16'd64919) begin
		isPrime = 1;
	end	else if (num==16'd64921) begin
		isPrime = 1;
	end	else if (num==16'd64927) begin
		isPrime = 1;
	end	else if (num==16'd64937) begin
		isPrime = 1;
	end	else if (num==16'd64951) begin
		isPrime = 1;
	end	else if (num==16'd64969) begin
		isPrime = 1;
	end	else if (num==16'd64997) begin
		isPrime = 1;
	end	else if (num==16'd65003) begin
		isPrime = 1;
	end	else if (num==16'd65011) begin
		isPrime = 1;
	end	else if (num==16'd65027) begin
		isPrime = 1;
	end	else if (num==16'd65029) begin
		isPrime = 1;
	end	else if (num==16'd65033) begin
		isPrime = 1;
	end	else if (num==16'd65053) begin
		isPrime = 1;
	end	else if (num==16'd65063) begin
		isPrime = 1;
	end	else if (num==16'd65071) begin
		isPrime = 1;
	end	else if (num==16'd65089) begin
		isPrime = 1;
	end	else if (num==16'd65099) begin
		isPrime = 1;
	end	else if (num==16'd65101) begin
		isPrime = 1;
	end	else if (num==16'd65111) begin
		isPrime = 1;
	end	else if (num==16'd65119) begin
		isPrime = 1;
	end	else if (num==16'd65123) begin
		isPrime = 1;
	end	else if (num==16'd65129) begin
		isPrime = 1;
	end	else if (num==16'd65141) begin
		isPrime = 1;
	end	else if (num==16'd65147) begin
		isPrime = 1;
	end	else if (num==16'd65167) begin
		isPrime = 1;
	end	else if (num==16'd65171) begin
		isPrime = 1;
	end	else if (num==16'd65173) begin
		isPrime = 1;
	end	else if (num==16'd65179) begin
		isPrime = 1;
	end	else if (num==16'd65183) begin
		isPrime = 1;
	end	else if (num==16'd65203) begin
		isPrime = 1;
	end	else if (num==16'd65213) begin
		isPrime = 1;
	end	else if (num==16'd65239) begin
		isPrime = 1;
	end	else if (num==16'd65257) begin
		isPrime = 1;
	end	else if (num==16'd65267) begin
		isPrime = 1;
	end	else if (num==16'd65269) begin
		isPrime = 1;
	end	else if (num==16'd65287) begin
		isPrime = 1;
	end	else if (num==16'd65293) begin
		isPrime = 1;
	end	else if (num==16'd65309) begin
		isPrime = 1;
	end	else if (num==16'd65323) begin
		isPrime = 1;
	end	else if (num==16'd65327) begin
		isPrime = 1;
	end	else if (num==16'd65353) begin
		isPrime = 1;
	end	else if (num==16'd65357) begin
		isPrime = 1;
	end	else if (num==16'd65371) begin
		isPrime = 1;
	end	else if (num==16'd65381) begin
		isPrime = 1;
	end	else if (num==16'd65393) begin
		isPrime = 1;
	end	else if (num==16'd65407) begin
		isPrime = 1;
	end	else if (num==16'd65413) begin
		isPrime = 1;
	end	else if (num==16'd65419) begin
		isPrime = 1;
	end	else if (num==16'd65423) begin
		isPrime = 1;
	end	else if (num==16'd65437) begin
		isPrime = 1;
	end	else if (num==16'd65447) begin
		isPrime = 1;
	end	else if (num==16'd65449) begin
		isPrime = 1;
	end	else if (num==16'd65479) begin
		isPrime = 1;
	end	else if (num==16'd65497) begin
		isPrime = 1;
	end	else if (num==16'd65519) begin
		isPrime = 1;
	end	else if (num==16'd65521) begin
		isPrime = 1;
	end
end


endmodule