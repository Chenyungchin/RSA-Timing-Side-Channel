module CheckPrime #(parameter WIDTH = 8) (
    // input
    input                    clk,
    input                    rst_n,
    input                    start,
    input      [  WIDTH-1:0] num,
    // output
    output reg               IsPrime,
    output reg               finish,
    output reg               AssumePrime
);

// there is 6542 primes < 65536
parameter PRIME_COUNT = 6542;

// stores the prime numbers that are smaller than 65536
parameter [0: 16*PRIME_COUNT-1] PrimeArray = {
    16'd2,
    16'd3,
    16'd5,
    16'd7,
    16'd11,
    16'd13,
    16'd17,
    16'd19,
    16'd23,
    16'd29,
    16'd31,
    16'd37,
    16'd41,
    16'd43,
    16'd47,
    16'd53,
    16'd59,
    16'd61,
    16'd67,
    16'd71,
    16'd73,
    16'd79,
    16'd83,
    16'd89,
    16'd97,
    16'd101,
    16'd103,
    16'd107,
    16'd109,
    16'd113,
    16'd127,
    16'd131,
    16'd137,
    16'd139,
    16'd149,
    16'd151,
    16'd157,
    16'd163,
    16'd167,
    16'd173,
    16'd179,
    16'd181,
    16'd191,
    16'd193,
    16'd197,
    16'd199,
    16'd211,
    16'd223,
    16'd227,
    16'd229,
    16'd233,
    16'd239,
    16'd241,
    16'd251,
    16'd257,
    16'd263,
    16'd269,
    16'd271,
    16'd277,
    16'd281,
    16'd283,
    16'd293,
    16'd307,
    16'd311,
    16'd313,
    16'd317,
    16'd331,
    16'd337,
    16'd347,
    16'd349,
    16'd353,
    16'd359,
    16'd367,
    16'd373,
    16'd379,
    16'd383,
    16'd389,
    16'd397,
    16'd401,
    16'd409,
    16'd419,
    16'd421,
    16'd431,
    16'd433,
    16'd439,
    16'd443,
    16'd449,
    16'd457,
    16'd461,
    16'd463,
    16'd467,
    16'd479,
    16'd487,
    16'd491,
    16'd499,
    16'd503,
    16'd509,
    16'd521,
    16'd523,
    16'd541,
    16'd547,
    16'd557,
    16'd563,
    16'd569,
    16'd571,
    16'd577,
    16'd587,
    16'd593,
    16'd599,
    16'd601,
    16'd607,
    16'd613,
    16'd617,
    16'd619,
    16'd631,
    16'd641,
    16'd643,
    16'd647,
    16'd653,
    16'd659,
    16'd661,
    16'd673,
    16'd677,
    16'd683,
    16'd691,
    16'd701,
    16'd709,
    16'd719,
    16'd727,
    16'd733,
    16'd739,
    16'd743,
    16'd751,
    16'd757,
    16'd761,
    16'd769,
    16'd773,
    16'd787,
    16'd797,
    16'd809,
    16'd811,
    16'd821,
    16'd823,
    16'd827,
    16'd829,
    16'd839,
    16'd853,
    16'd857,
    16'd859,
    16'd863,
    16'd877,
    16'd881,
    16'd883,
    16'd887,
    16'd907,
    16'd911,
    16'd919,
    16'd929,
    16'd937,
    16'd941,
    16'd947,
    16'd953,
    16'd967,
    16'd971,
    16'd977,
    16'd983,
    16'd991,
    16'd997,
    16'd1009,
    16'd1013,
    16'd1019,
    16'd1021,
    16'd1031,
    16'd1033,
    16'd1039,
    16'd1049,
    16'd1051,
    16'd1061,
    16'd1063,
    16'd1069,
    16'd1087,
    16'd1091,
    16'd1093,
    16'd1097,
    16'd1103,
    16'd1109,
    16'd1117,
    16'd1123,
    16'd1129,
    16'd1151,
    16'd1153,
    16'd1163,
    16'd1171,
    16'd1181,
    16'd1187,
    16'd1193,
    16'd1201,
    16'd1213,
    16'd1217,
    16'd1223,
    16'd1229,
    16'd1231,
    16'd1237,
    16'd1249,
    16'd1259,
    16'd1277,
    16'd1279,
    16'd1283,
    16'd1289,
    16'd1291,
    16'd1297,
    16'd1301,
    16'd1303,
    16'd1307,
    16'd1319,
    16'd1321,
    16'd1327,
    16'd1361,
    16'd1367,
    16'd1373,
    16'd1381,
    16'd1399,
    16'd1409,
    16'd1423,
    16'd1427,
    16'd1429,
    16'd1433,
    16'd1439,
    16'd1447,
    16'd1451,
    16'd1453,
    16'd1459,
    16'd1471,
    16'd1481,
    16'd1483,
    16'd1487,
    16'd1489,
    16'd1493,
    16'd1499,
    16'd1511,
    16'd1523,
    16'd1531,
    16'd1543,
    16'd1549,
    16'd1553,
    16'd1559,
    16'd1567,
    16'd1571,
    16'd1579,
    16'd1583,
    16'd1597,
    16'd1601,
    16'd1607,
    16'd1609,
    16'd1613,
    16'd1619,
    16'd1621,
    16'd1627,
    16'd1637,
    16'd1657,
    16'd1663,
    16'd1667,
    16'd1669,
    16'd1693,
    16'd1697,
    16'd1699,
    16'd1709,
    16'd1721,
    16'd1723,
    16'd1733,
    16'd1741,
    16'd1747,
    16'd1753,
    16'd1759,
    16'd1777,
    16'd1783,
    16'd1787,
    16'd1789,
    16'd1801,
    16'd1811,
    16'd1823,
    16'd1831,
    16'd1847,
    16'd1861,
    16'd1867,
    16'd1871,
    16'd1873,
    16'd1877,
    16'd1879,
    16'd1889,
    16'd1901,
    16'd1907,
    16'd1913,
    16'd1931,
    16'd1933,
    16'd1949,
    16'd1951,
    16'd1973,
    16'd1979,
    16'd1987,
    16'd1993,
    16'd1997,
    16'd1999,
    16'd2003,
    16'd2011,
    16'd2017,
    16'd2027,
    16'd2029,
    16'd2039,
    16'd2053,
    16'd2063,
    16'd2069,
    16'd2081,
    16'd2083,
    16'd2087,
    16'd2089,
    16'd2099,
    16'd2111,
    16'd2113,
    16'd2129,
    16'd2131,
    16'd2137,
    16'd2141,
    16'd2143,
    16'd2153,
    16'd2161,
    16'd2179,
    16'd2203,
    16'd2207,
    16'd2213,
    16'd2221,
    16'd2237,
    16'd2239,
    16'd2243,
    16'd2251,
    16'd2267,
    16'd2269,
    16'd2273,
    16'd2281,
    16'd2287,
    16'd2293,
    16'd2297,
    16'd2309,
    16'd2311,
    16'd2333,
    16'd2339,
    16'd2341,
    16'd2347,
    16'd2351,
    16'd2357,
    16'd2371,
    16'd2377,
    16'd2381,
    16'd2383,
    16'd2389,
    16'd2393,
    16'd2399,
    16'd2411,
    16'd2417,
    16'd2423,
    16'd2437,
    16'd2441,
    16'd2447,
    16'd2459,
    16'd2467,
    16'd2473,
    16'd2477,
    16'd2503,
    16'd2521,
    16'd2531,
    16'd2539,
    16'd2543,
    16'd2549,
    16'd2551,
    16'd2557,
    16'd2579,
    16'd2591,
    16'd2593,
    16'd2609,
    16'd2617,
    16'd2621,
    16'd2633,
    16'd2647,
    16'd2657,
    16'd2659,
    16'd2663,
    16'd2671,
    16'd2677,
    16'd2683,
    16'd2687,
    16'd2689,
    16'd2693,
    16'd2699,
    16'd2707,
    16'd2711,
    16'd2713,
    16'd2719,
    16'd2729,
    16'd2731,
    16'd2741,
    16'd2749,
    16'd2753,
    16'd2767,
    16'd2777,
    16'd2789,
    16'd2791,
    16'd2797,
    16'd2801,
    16'd2803,
    16'd2819,
    16'd2833,
    16'd2837,
    16'd2843,
    16'd2851,
    16'd2857,
    16'd2861,
    16'd2879,
    16'd2887,
    16'd2897,
    16'd2903,
    16'd2909,
    16'd2917,
    16'd2927,
    16'd2939,
    16'd2953,
    16'd2957,
    16'd2963,
    16'd2969,
    16'd2971,
    16'd2999,
    16'd3001,
    16'd3011,
    16'd3019,
    16'd3023,
    16'd3037,
    16'd3041,
    16'd3049,
    16'd3061,
    16'd3067,
    16'd3079,
    16'd3083,
    16'd3089,
    16'd3109,
    16'd3119,
    16'd3121,
    16'd3137,
    16'd3163,
    16'd3167,
    16'd3169,
    16'd3181,
    16'd3187,
    16'd3191,
    16'd3203,
    16'd3209,
    16'd3217,
    16'd3221,
    16'd3229,
    16'd3251,
    16'd3253,
    16'd3257,
    16'd3259,
    16'd3271,
    16'd3299,
    16'd3301,
    16'd3307,
    16'd3313,
    16'd3319,
    16'd3323,
    16'd3329,
    16'd3331,
    16'd3343,
    16'd3347,
    16'd3359,
    16'd3361,
    16'd3371,
    16'd3373,
    16'd3389,
    16'd3391,
    16'd3407,
    16'd3413,
    16'd3433,
    16'd3449,
    16'd3457,
    16'd3461,
    16'd3463,
    16'd3467,
    16'd3469,
    16'd3491,
    16'd3499,
    16'd3511,
    16'd3517,
    16'd3527,
    16'd3529,
    16'd3533,
    16'd3539,
    16'd3541,
    16'd3547,
    16'd3557,
    16'd3559,
    16'd3571,
    16'd3581,
    16'd3583,
    16'd3593,
    16'd3607,
    16'd3613,
    16'd3617,
    16'd3623,
    16'd3631,
    16'd3637,
    16'd3643,
    16'd3659,
    16'd3671,
    16'd3673,
    16'd3677,
    16'd3691,
    16'd3697,
    16'd3701,
    16'd3709,
    16'd3719,
    16'd3727,
    16'd3733,
    16'd3739,
    16'd3761,
    16'd3767,
    16'd3769,
    16'd3779,
    16'd3793,
    16'd3797,
    16'd3803,
    16'd3821,
    16'd3823,
    16'd3833,
    16'd3847,
    16'd3851,
    16'd3853,
    16'd3863,
    16'd3877,
    16'd3881,
    16'd3889,
    16'd3907,
    16'd3911,
    16'd3917,
    16'd3919,
    16'd3923,
    16'd3929,
    16'd3931,
    16'd3943,
    16'd3947,
    16'd3967,
    16'd3989,
    16'd4001,
    16'd4003,
    16'd4007,
    16'd4013,
    16'd4019,
    16'd4021,
    16'd4027,
    16'd4049,
    16'd4051,
    16'd4057,
    16'd4073,
    16'd4079,
    16'd4091,
    16'd4093,
    16'd4099,
    16'd4111,
    16'd4127,
    16'd4129,
    16'd4133,
    16'd4139,
    16'd4153,
    16'd4157,
    16'd4159,
    16'd4177,
    16'd4201,
    16'd4211,
    16'd4217,
    16'd4219,
    16'd4229,
    16'd4231,
    16'd4241,
    16'd4243,
    16'd4253,
    16'd4259,
    16'd4261,
    16'd4271,
    16'd4273,
    16'd4283,
    16'd4289,
    16'd4297,
    16'd4327,
    16'd4337,
    16'd4339,
    16'd4349,
    16'd4357,
    16'd4363,
    16'd4373,
    16'd4391,
    16'd4397,
    16'd4409,
    16'd4421,
    16'd4423,
    16'd4441,
    16'd4447,
    16'd4451,
    16'd4457,
    16'd4463,
    16'd4481,
    16'd4483,
    16'd4493,
    16'd4507,
    16'd4513,
    16'd4517,
    16'd4519,
    16'd4523,
    16'd4547,
    16'd4549,
    16'd4561,
    16'd4567,
    16'd4583,
    16'd4591,
    16'd4597,
    16'd4603,
    16'd4621,
    16'd4637,
    16'd4639,
    16'd4643,
    16'd4649,
    16'd4651,
    16'd4657,
    16'd4663,
    16'd4673,
    16'd4679,
    16'd4691,
    16'd4703,
    16'd4721,
    16'd4723,
    16'd4729,
    16'd4733,
    16'd4751,
    16'd4759,
    16'd4783,
    16'd4787,
    16'd4789,
    16'd4793,
    16'd4799,
    16'd4801,
    16'd4813,
    16'd4817,
    16'd4831,
    16'd4861,
    16'd4871,
    16'd4877,
    16'd4889,
    16'd4903,
    16'd4909,
    16'd4919,
    16'd4931,
    16'd4933,
    16'd4937,
    16'd4943,
    16'd4951,
    16'd4957,
    16'd4967,
    16'd4969,
    16'd4973,
    16'd4987,
    16'd4993,
    16'd4999,
    16'd5003,
    16'd5009,
    16'd5011,
    16'd5021,
    16'd5023,
    16'd5039,
    16'd5051,
    16'd5059,
    16'd5077,
    16'd5081,
    16'd5087,
    16'd5099,
    16'd5101,
    16'd5107,
    16'd5113,
    16'd5119,
    16'd5147,
    16'd5153,
    16'd5167,
    16'd5171,
    16'd5179,
    16'd5189,
    16'd5197,
    16'd5209,
    16'd5227,
    16'd5231,
    16'd5233,
    16'd5237,
    16'd5261,
    16'd5273,
    16'd5279,
    16'd5281,
    16'd5297,
    16'd5303,
    16'd5309,
    16'd5323,
    16'd5333,
    16'd5347,
    16'd5351,
    16'd5381,
    16'd5387,
    16'd5393,
    16'd5399,
    16'd5407,
    16'd5413,
    16'd5417,
    16'd5419,
    16'd5431,
    16'd5437,
    16'd5441,
    16'd5443,
    16'd5449,
    16'd5471,
    16'd5477,
    16'd5479,
    16'd5483,
    16'd5501,
    16'd5503,
    16'd5507,
    16'd5519,
    16'd5521,
    16'd5527,
    16'd5531,
    16'd5557,
    16'd5563,
    16'd5569,
    16'd5573,
    16'd5581,
    16'd5591,
    16'd5623,
    16'd5639,
    16'd5641,
    16'd5647,
    16'd5651,
    16'd5653,
    16'd5657,
    16'd5659,
    16'd5669,
    16'd5683,
    16'd5689,
    16'd5693,
    16'd5701,
    16'd5711,
    16'd5717,
    16'd5737,
    16'd5741,
    16'd5743,
    16'd5749,
    16'd5779,
    16'd5783,
    16'd5791,
    16'd5801,
    16'd5807,
    16'd5813,
    16'd5821,
    16'd5827,
    16'd5839,
    16'd5843,
    16'd5849,
    16'd5851,
    16'd5857,
    16'd5861,
    16'd5867,
    16'd5869,
    16'd5879,
    16'd5881,
    16'd5897,
    16'd5903,
    16'd5923,
    16'd5927,
    16'd5939,
    16'd5953,
    16'd5981,
    16'd5987,
    16'd6007,
    16'd6011,
    16'd6029,
    16'd6037,
    16'd6043,
    16'd6047,
    16'd6053,
    16'd6067,
    16'd6073,
    16'd6079,
    16'd6089,
    16'd6091,
    16'd6101,
    16'd6113,
    16'd6121,
    16'd6131,
    16'd6133,
    16'd6143,
    16'd6151,
    16'd6163,
    16'd6173,
    16'd6197,
    16'd6199,
    16'd6203,
    16'd6211,
    16'd6217,
    16'd6221,
    16'd6229,
    16'd6247,
    16'd6257,
    16'd6263,
    16'd6269,
    16'd6271,
    16'd6277,
    16'd6287,
    16'd6299,
    16'd6301,
    16'd6311,
    16'd6317,
    16'd6323,
    16'd6329,
    16'd6337,
    16'd6343,
    16'd6353,
    16'd6359,
    16'd6361,
    16'd6367,
    16'd6373,
    16'd6379,
    16'd6389,
    16'd6397,
    16'd6421,
    16'd6427,
    16'd6449,
    16'd6451,
    16'd6469,
    16'd6473,
    16'd6481,
    16'd6491,
    16'd6521,
    16'd6529,
    16'd6547,
    16'd6551,
    16'd6553,
    16'd6563,
    16'd6569,
    16'd6571,
    16'd6577,
    16'd6581,
    16'd6599,
    16'd6607,
    16'd6619,
    16'd6637,
    16'd6653,
    16'd6659,
    16'd6661,
    16'd6673,
    16'd6679,
    16'd6689,
    16'd6691,
    16'd6701,
    16'd6703,
    16'd6709,
    16'd6719,
    16'd6733,
    16'd6737,
    16'd6761,
    16'd6763,
    16'd6779,
    16'd6781,
    16'd6791,
    16'd6793,
    16'd6803,
    16'd6823,
    16'd6827,
    16'd6829,
    16'd6833,
    16'd6841,
    16'd6857,
    16'd6863,
    16'd6869,
    16'd6871,
    16'd6883,
    16'd6899,
    16'd6907,
    16'd6911,
    16'd6917,
    16'd6947,
    16'd6949,
    16'd6959,
    16'd6961,
    16'd6967,
    16'd6971,
    16'd6977,
    16'd6983,
    16'd6991,
    16'd6997,
    16'd7001,
    16'd7013,
    16'd7019,
    16'd7027,
    16'd7039,
    16'd7043,
    16'd7057,
    16'd7069,
    16'd7079,
    16'd7103,
    16'd7109,
    16'd7121,
    16'd7127,
    16'd7129,
    16'd7151,
    16'd7159,
    16'd7177,
    16'd7187,
    16'd7193,
    16'd7207,
    16'd7211,
    16'd7213,
    16'd7219,
    16'd7229,
    16'd7237,
    16'd7243,
    16'd7247,
    16'd7253,
    16'd7283,
    16'd7297,
    16'd7307,
    16'd7309,
    16'd7321,
    16'd7331,
    16'd7333,
    16'd7349,
    16'd7351,
    16'd7369,
    16'd7393,
    16'd7411,
    16'd7417,
    16'd7433,
    16'd7451,
    16'd7457,
    16'd7459,
    16'd7477,
    16'd7481,
    16'd7487,
    16'd7489,
    16'd7499,
    16'd7507,
    16'd7517,
    16'd7523,
    16'd7529,
    16'd7537,
    16'd7541,
    16'd7547,
    16'd7549,
    16'd7559,
    16'd7561,
    16'd7573,
    16'd7577,
    16'd7583,
    16'd7589,
    16'd7591,
    16'd7603,
    16'd7607,
    16'd7621,
    16'd7639,
    16'd7643,
    16'd7649,
    16'd7669,
    16'd7673,
    16'd7681,
    16'd7687,
    16'd7691,
    16'd7699,
    16'd7703,
    16'd7717,
    16'd7723,
    16'd7727,
    16'd7741,
    16'd7753,
    16'd7757,
    16'd7759,
    16'd7789,
    16'd7793,
    16'd7817,
    16'd7823,
    16'd7829,
    16'd7841,
    16'd7853,
    16'd7867,
    16'd7873,
    16'd7877,
    16'd7879,
    16'd7883,
    16'd7901,
    16'd7907,
    16'd7919,
    16'd7927,
    16'd7933,
    16'd7937,
    16'd7949,
    16'd7951,
    16'd7963,
    16'd7993,
    16'd8009,
    16'd8011,
    16'd8017,
    16'd8039,
    16'd8053,
    16'd8059,
    16'd8069,
    16'd8081,
    16'd8087,
    16'd8089,
    16'd8093,
    16'd8101,
    16'd8111,
    16'd8117,
    16'd8123,
    16'd8147,
    16'd8161,
    16'd8167,
    16'd8171,
    16'd8179,
    16'd8191,
    16'd8209,
    16'd8219,
    16'd8221,
    16'd8231,
    16'd8233,
    16'd8237,
    16'd8243,
    16'd8263,
    16'd8269,
    16'd8273,
    16'd8287,
    16'd8291,
    16'd8293,
    16'd8297,
    16'd8311,
    16'd8317,
    16'd8329,
    16'd8353,
    16'd8363,
    16'd8369,
    16'd8377,
    16'd8387,
    16'd8389,
    16'd8419,
    16'd8423,
    16'd8429,
    16'd8431,
    16'd8443,
    16'd8447,
    16'd8461,
    16'd8467,
    16'd8501,
    16'd8513,
    16'd8521,
    16'd8527,
    16'd8537,
    16'd8539,
    16'd8543,
    16'd8563,
    16'd8573,
    16'd8581,
    16'd8597,
    16'd8599,
    16'd8609,
    16'd8623,
    16'd8627,
    16'd8629,
    16'd8641,
    16'd8647,
    16'd8663,
    16'd8669,
    16'd8677,
    16'd8681,
    16'd8689,
    16'd8693,
    16'd8699,
    16'd8707,
    16'd8713,
    16'd8719,
    16'd8731,
    16'd8737,
    16'd8741,
    16'd8747,
    16'd8753,
    16'd8761,
    16'd8779,
    16'd8783,
    16'd8803,
    16'd8807,
    16'd8819,
    16'd8821,
    16'd8831,
    16'd8837,
    16'd8839,
    16'd8849,
    16'd8861,
    16'd8863,
    16'd8867,
    16'd8887,
    16'd8893,
    16'd8923,
    16'd8929,
    16'd8933,
    16'd8941,
    16'd8951,
    16'd8963,
    16'd8969,
    16'd8971,
    16'd8999,
    16'd9001,
    16'd9007,
    16'd9011,
    16'd9013,
    16'd9029,
    16'd9041,
    16'd9043,
    16'd9049,
    16'd9059,
    16'd9067,
    16'd9091,
    16'd9103,
    16'd9109,
    16'd9127,
    16'd9133,
    16'd9137,
    16'd9151,
    16'd9157,
    16'd9161,
    16'd9173,
    16'd9181,
    16'd9187,
    16'd9199,
    16'd9203,
    16'd9209,
    16'd9221,
    16'd9227,
    16'd9239,
    16'd9241,
    16'd9257,
    16'd9277,
    16'd9281,
    16'd9283,
    16'd9293,
    16'd9311,
    16'd9319,
    16'd9323,
    16'd9337,
    16'd9341,
    16'd9343,
    16'd9349,
    16'd9371,
    16'd9377,
    16'd9391,
    16'd9397,
    16'd9403,
    16'd9413,
    16'd9419,
    16'd9421,
    16'd9431,
    16'd9433,
    16'd9437,
    16'd9439,
    16'd9461,
    16'd9463,
    16'd9467,
    16'd9473,
    16'd9479,
    16'd9491,
    16'd9497,
    16'd9511,
    16'd9521,
    16'd9533,
    16'd9539,
    16'd9547,
    16'd9551,
    16'd9587,
    16'd9601,
    16'd9613,
    16'd9619,
    16'd9623,
    16'd9629,
    16'd9631,
    16'd9643,
    16'd9649,
    16'd9661,
    16'd9677,
    16'd9679,
    16'd9689,
    16'd9697,
    16'd9719,
    16'd9721,
    16'd9733,
    16'd9739,
    16'd9743,
    16'd9749,
    16'd9767,
    16'd9769,
    16'd9781,
    16'd9787,
    16'd9791,
    16'd9803,
    16'd9811,
    16'd9817,
    16'd9829,
    16'd9833,
    16'd9839,
    16'd9851,
    16'd9857,
    16'd9859,
    16'd9871,
    16'd9883,
    16'd9887,
    16'd9901,
    16'd9907,
    16'd9923,
    16'd9929,
    16'd9931,
    16'd9941,
    16'd9949,
    16'd9967,
    16'd9973,
    16'd10007,
    16'd10009,
    16'd10037,
    16'd10039,
    16'd10061,
    16'd10067,
    16'd10069,
    16'd10079,
    16'd10091,
    16'd10093,
    16'd10099,
    16'd10103,
    16'd10111,
    16'd10133,
    16'd10139,
    16'd10141,
    16'd10151,
    16'd10159,
    16'd10163,
    16'd10169,
    16'd10177,
    16'd10181,
    16'd10193,
    16'd10211,
    16'd10223,
    16'd10243,
    16'd10247,
    16'd10253,
    16'd10259,
    16'd10267,
    16'd10271,
    16'd10273,
    16'd10289,
    16'd10301,
    16'd10303,
    16'd10313,
    16'd10321,
    16'd10331,
    16'd10333,
    16'd10337,
    16'd10343,
    16'd10357,
    16'd10369,
    16'd10391,
    16'd10399,
    16'd10427,
    16'd10429,
    16'd10433,
    16'd10453,
    16'd10457,
    16'd10459,
    16'd10463,
    16'd10477,
    16'd10487,
    16'd10499,
    16'd10501,
    16'd10513,
    16'd10529,
    16'd10531,
    16'd10559,
    16'd10567,
    16'd10589,
    16'd10597,
    16'd10601,
    16'd10607,
    16'd10613,
    16'd10627,
    16'd10631,
    16'd10639,
    16'd10651,
    16'd10657,
    16'd10663,
    16'd10667,
    16'd10687,
    16'd10691,
    16'd10709,
    16'd10711,
    16'd10723,
    16'd10729,
    16'd10733,
    16'd10739,
    16'd10753,
    16'd10771,
    16'd10781,
    16'd10789,
    16'd10799,
    16'd10831,
    16'd10837,
    16'd10847,
    16'd10853,
    16'd10859,
    16'd10861,
    16'd10867,
    16'd10883,
    16'd10889,
    16'd10891,
    16'd10903,
    16'd10909,
    16'd10937,
    16'd10939,
    16'd10949,
    16'd10957,
    16'd10973,
    16'd10979,
    16'd10987,
    16'd10993,
    16'd11003,
    16'd11027,
    16'd11047,
    16'd11057,
    16'd11059,
    16'd11069,
    16'd11071,
    16'd11083,
    16'd11087,
    16'd11093,
    16'd11113,
    16'd11117,
    16'd11119,
    16'd11131,
    16'd11149,
    16'd11159,
    16'd11161,
    16'd11171,
    16'd11173,
    16'd11177,
    16'd11197,
    16'd11213,
    16'd11239,
    16'd11243,
    16'd11251,
    16'd11257,
    16'd11261,
    16'd11273,
    16'd11279,
    16'd11287,
    16'd11299,
    16'd11311,
    16'd11317,
    16'd11321,
    16'd11329,
    16'd11351,
    16'd11353,
    16'd11369,
    16'd11383,
    16'd11393,
    16'd11399,
    16'd11411,
    16'd11423,
    16'd11437,
    16'd11443,
    16'd11447,
    16'd11467,
    16'd11471,
    16'd11483,
    16'd11489,
    16'd11491,
    16'd11497,
    16'd11503,
    16'd11519,
    16'd11527,
    16'd11549,
    16'd11551,
    16'd11579,
    16'd11587,
    16'd11593,
    16'd11597,
    16'd11617,
    16'd11621,
    16'd11633,
    16'd11657,
    16'd11677,
    16'd11681,
    16'd11689,
    16'd11699,
    16'd11701,
    16'd11717,
    16'd11719,
    16'd11731,
    16'd11743,
    16'd11777,
    16'd11779,
    16'd11783,
    16'd11789,
    16'd11801,
    16'd11807,
    16'd11813,
    16'd11821,
    16'd11827,
    16'd11831,
    16'd11833,
    16'd11839,
    16'd11863,
    16'd11867,
    16'd11887,
    16'd11897,
    16'd11903,
    16'd11909,
    16'd11923,
    16'd11927,
    16'd11933,
    16'd11939,
    16'd11941,
    16'd11953,
    16'd11959,
    16'd11969,
    16'd11971,
    16'd11981,
    16'd11987,
    16'd12007,
    16'd12011,
    16'd12037,
    16'd12041,
    16'd12043,
    16'd12049,
    16'd12071,
    16'd12073,
    16'd12097,
    16'd12101,
    16'd12107,
    16'd12109,
    16'd12113,
    16'd12119,
    16'd12143,
    16'd12149,
    16'd12157,
    16'd12161,
    16'd12163,
    16'd12197,
    16'd12203,
    16'd12211,
    16'd12227,
    16'd12239,
    16'd12241,
    16'd12251,
    16'd12253,
    16'd12263,
    16'd12269,
    16'd12277,
    16'd12281,
    16'd12289,
    16'd12301,
    16'd12323,
    16'd12329,
    16'd12343,
    16'd12347,
    16'd12373,
    16'd12377,
    16'd12379,
    16'd12391,
    16'd12401,
    16'd12409,
    16'd12413,
    16'd12421,
    16'd12433,
    16'd12437,
    16'd12451,
    16'd12457,
    16'd12473,
    16'd12479,
    16'd12487,
    16'd12491,
    16'd12497,
    16'd12503,
    16'd12511,
    16'd12517,
    16'd12527,
    16'd12539,
    16'd12541,
    16'd12547,
    16'd12553,
    16'd12569,
    16'd12577,
    16'd12583,
    16'd12589,
    16'd12601,
    16'd12611,
    16'd12613,
    16'd12619,
    16'd12637,
    16'd12641,
    16'd12647,
    16'd12653,
    16'd12659,
    16'd12671,
    16'd12689,
    16'd12697,
    16'd12703,
    16'd12713,
    16'd12721,
    16'd12739,
    16'd12743,
    16'd12757,
    16'd12763,
    16'd12781,
    16'd12791,
    16'd12799,
    16'd12809,
    16'd12821,
    16'd12823,
    16'd12829,
    16'd12841,
    16'd12853,
    16'd12889,
    16'd12893,
    16'd12899,
    16'd12907,
    16'd12911,
    16'd12917,
    16'd12919,
    16'd12923,
    16'd12941,
    16'd12953,
    16'd12959,
    16'd12967,
    16'd12973,
    16'd12979,
    16'd12983,
    16'd13001,
    16'd13003,
    16'd13007,
    16'd13009,
    16'd13033,
    16'd13037,
    16'd13043,
    16'd13049,
    16'd13063,
    16'd13093,
    16'd13099,
    16'd13103,
    16'd13109,
    16'd13121,
    16'd13127,
    16'd13147,
    16'd13151,
    16'd13159,
    16'd13163,
    16'd13171,
    16'd13177,
    16'd13183,
    16'd13187,
    16'd13217,
    16'd13219,
    16'd13229,
    16'd13241,
    16'd13249,
    16'd13259,
    16'd13267,
    16'd13291,
    16'd13297,
    16'd13309,
    16'd13313,
    16'd13327,
    16'd13331,
    16'd13337,
    16'd13339,
    16'd13367,
    16'd13381,
    16'd13397,
    16'd13399,
    16'd13411,
    16'd13417,
    16'd13421,
    16'd13441,
    16'd13451,
    16'd13457,
    16'd13463,
    16'd13469,
    16'd13477,
    16'd13487,
    16'd13499,
    16'd13513,
    16'd13523,
    16'd13537,
    16'd13553,
    16'd13567,
    16'd13577,
    16'd13591,
    16'd13597,
    16'd13613,
    16'd13619,
    16'd13627,
    16'd13633,
    16'd13649,
    16'd13669,
    16'd13679,
    16'd13681,
    16'd13687,
    16'd13691,
    16'd13693,
    16'd13697,
    16'd13709,
    16'd13711,
    16'd13721,
    16'd13723,
    16'd13729,
    16'd13751,
    16'd13757,
    16'd13759,
    16'd13763,
    16'd13781,
    16'd13789,
    16'd13799,
    16'd13807,
    16'd13829,
    16'd13831,
    16'd13841,
    16'd13859,
    16'd13873,
    16'd13877,
    16'd13879,
    16'd13883,
    16'd13901,
    16'd13903,
    16'd13907,
    16'd13913,
    16'd13921,
    16'd13931,
    16'd13933,
    16'd13963,
    16'd13967,
    16'd13997,
    16'd13999,
    16'd14009,
    16'd14011,
    16'd14029,
    16'd14033,
    16'd14051,
    16'd14057,
    16'd14071,
    16'd14081,
    16'd14083,
    16'd14087,
    16'd14107,
    16'd14143,
    16'd14149,
    16'd14153,
    16'd14159,
    16'd14173,
    16'd14177,
    16'd14197,
    16'd14207,
    16'd14221,
    16'd14243,
    16'd14249,
    16'd14251,
    16'd14281,
    16'd14293,
    16'd14303,
    16'd14321,
    16'd14323,
    16'd14327,
    16'd14341,
    16'd14347,
    16'd14369,
    16'd14387,
    16'd14389,
    16'd14401,
    16'd14407,
    16'd14411,
    16'd14419,
    16'd14423,
    16'd14431,
    16'd14437,
    16'd14447,
    16'd14449,
    16'd14461,
    16'd14479,
    16'd14489,
    16'd14503,
    16'd14519,
    16'd14533,
    16'd14537,
    16'd14543,
    16'd14549,
    16'd14551,
    16'd14557,
    16'd14561,
    16'd14563,
    16'd14591,
    16'd14593,
    16'd14621,
    16'd14627,
    16'd14629,
    16'd14633,
    16'd14639,
    16'd14653,
    16'd14657,
    16'd14669,
    16'd14683,
    16'd14699,
    16'd14713,
    16'd14717,
    16'd14723,
    16'd14731,
    16'd14737,
    16'd14741,
    16'd14747,
    16'd14753,
    16'd14759,
    16'd14767,
    16'd14771,
    16'd14779,
    16'd14783,
    16'd14797,
    16'd14813,
    16'd14821,
    16'd14827,
    16'd14831,
    16'd14843,
    16'd14851,
    16'd14867,
    16'd14869,
    16'd14879,
    16'd14887,
    16'd14891,
    16'd14897,
    16'd14923,
    16'd14929,
    16'd14939,
    16'd14947,
    16'd14951,
    16'd14957,
    16'd14969,
    16'd14983,
    16'd15013,
    16'd15017,
    16'd15031,
    16'd15053,
    16'd15061,
    16'd15073,
    16'd15077,
    16'd15083,
    16'd15091,
    16'd15101,
    16'd15107,
    16'd15121,
    16'd15131,
    16'd15137,
    16'd15139,
    16'd15149,
    16'd15161,
    16'd15173,
    16'd15187,
    16'd15193,
    16'd15199,
    16'd15217,
    16'd15227,
    16'd15233,
    16'd15241,
    16'd15259,
    16'd15263,
    16'd15269,
    16'd15271,
    16'd15277,
    16'd15287,
    16'd15289,
    16'd15299,
    16'd15307,
    16'd15313,
    16'd15319,
    16'd15329,
    16'd15331,
    16'd15349,
    16'd15359,
    16'd15361,
    16'd15373,
    16'd15377,
    16'd15383,
    16'd15391,
    16'd15401,
    16'd15413,
    16'd15427,
    16'd15439,
    16'd15443,
    16'd15451,
    16'd15461,
    16'd15467,
    16'd15473,
    16'd15493,
    16'd15497,
    16'd15511,
    16'd15527,
    16'd15541,
    16'd15551,
    16'd15559,
    16'd15569,
    16'd15581,
    16'd15583,
    16'd15601,
    16'd15607,
    16'd15619,
    16'd15629,
    16'd15641,
    16'd15643,
    16'd15647,
    16'd15649,
    16'd15661,
    16'd15667,
    16'd15671,
    16'd15679,
    16'd15683,
    16'd15727,
    16'd15731,
    16'd15733,
    16'd15737,
    16'd15739,
    16'd15749,
    16'd15761,
    16'd15767,
    16'd15773,
    16'd15787,
    16'd15791,
    16'd15797,
    16'd15803,
    16'd15809,
    16'd15817,
    16'd15823,
    16'd15859,
    16'd15877,
    16'd15881,
    16'd15887,
    16'd15889,
    16'd15901,
    16'd15907,
    16'd15913,
    16'd15919,
    16'd15923,
    16'd15937,
    16'd15959,
    16'd15971,
    16'd15973,
    16'd15991,
    16'd16001,
    16'd16007,
    16'd16033,
    16'd16057,
    16'd16061,
    16'd16063,
    16'd16067,
    16'd16069,
    16'd16073,
    16'd16087,
    16'd16091,
    16'd16097,
    16'd16103,
    16'd16111,
    16'd16127,
    16'd16139,
    16'd16141,
    16'd16183,
    16'd16187,
    16'd16189,
    16'd16193,
    16'd16217,
    16'd16223,
    16'd16229,
    16'd16231,
    16'd16249,
    16'd16253,
    16'd16267,
    16'd16273,
    16'd16301,
    16'd16319,
    16'd16333,
    16'd16339,
    16'd16349,
    16'd16361,
    16'd16363,
    16'd16369,
    16'd16381,
    16'd16411,
    16'd16417,
    16'd16421,
    16'd16427,
    16'd16433,
    16'd16447,
    16'd16451,
    16'd16453,
    16'd16477,
    16'd16481,
    16'd16487,
    16'd16493,
    16'd16519,
    16'd16529,
    16'd16547,
    16'd16553,
    16'd16561,
    16'd16567,
    16'd16573,
    16'd16603,
    16'd16607,
    16'd16619,
    16'd16631,
    16'd16633,
    16'd16649,
    16'd16651,
    16'd16657,
    16'd16661,
    16'd16673,
    16'd16691,
    16'd16693,
    16'd16699,
    16'd16703,
    16'd16729,
    16'd16741,
    16'd16747,
    16'd16759,
    16'd16763,
    16'd16787,
    16'd16811,
    16'd16823,
    16'd16829,
    16'd16831,
    16'd16843,
    16'd16871,
    16'd16879,
    16'd16883,
    16'd16889,
    16'd16901,
    16'd16903,
    16'd16921,
    16'd16927,
    16'd16931,
    16'd16937,
    16'd16943,
    16'd16963,
    16'd16979,
    16'd16981,
    16'd16987,
    16'd16993,
    16'd17011,
    16'd17021,
    16'd17027,
    16'd17029,
    16'd17033,
    16'd17041,
    16'd17047,
    16'd17053,
    16'd17077,
    16'd17093,
    16'd17099,
    16'd17107,
    16'd17117,
    16'd17123,
    16'd17137,
    16'd17159,
    16'd17167,
    16'd17183,
    16'd17189,
    16'd17191,
    16'd17203,
    16'd17207,
    16'd17209,
    16'd17231,
    16'd17239,
    16'd17257,
    16'd17291,
    16'd17293,
    16'd17299,
    16'd17317,
    16'd17321,
    16'd17327,
    16'd17333,
    16'd17341,
    16'd17351,
    16'd17359,
    16'd17377,
    16'd17383,
    16'd17387,
    16'd17389,
    16'd17393,
    16'd17401,
    16'd17417,
    16'd17419,
    16'd17431,
    16'd17443,
    16'd17449,
    16'd17467,
    16'd17471,
    16'd17477,
    16'd17483,
    16'd17489,
    16'd17491,
    16'd17497,
    16'd17509,
    16'd17519,
    16'd17539,
    16'd17551,
    16'd17569,
    16'd17573,
    16'd17579,
    16'd17581,
    16'd17597,
    16'd17599,
    16'd17609,
    16'd17623,
    16'd17627,
    16'd17657,
    16'd17659,
    16'd17669,
    16'd17681,
    16'd17683,
    16'd17707,
    16'd17713,
    16'd17729,
    16'd17737,
    16'd17747,
    16'd17749,
    16'd17761,
    16'd17783,
    16'd17789,
    16'd17791,
    16'd17807,
    16'd17827,
    16'd17837,
    16'd17839,
    16'd17851,
    16'd17863,
    16'd17881,
    16'd17891,
    16'd17903,
    16'd17909,
    16'd17911,
    16'd17921,
    16'd17923,
    16'd17929,
    16'd17939,
    16'd17957,
    16'd17959,
    16'd17971,
    16'd17977,
    16'd17981,
    16'd17987,
    16'd17989,
    16'd18013,
    16'd18041,
    16'd18043,
    16'd18047,
    16'd18049,
    16'd18059,
    16'd18061,
    16'd18077,
    16'd18089,
    16'd18097,
    16'd18119,
    16'd18121,
    16'd18127,
    16'd18131,
    16'd18133,
    16'd18143,
    16'd18149,
    16'd18169,
    16'd18181,
    16'd18191,
    16'd18199,
    16'd18211,
    16'd18217,
    16'd18223,
    16'd18229,
    16'd18233,
    16'd18251,
    16'd18253,
    16'd18257,
    16'd18269,
    16'd18287,
    16'd18289,
    16'd18301,
    16'd18307,
    16'd18311,
    16'd18313,
    16'd18329,
    16'd18341,
    16'd18353,
    16'd18367,
    16'd18371,
    16'd18379,
    16'd18397,
    16'd18401,
    16'd18413,
    16'd18427,
    16'd18433,
    16'd18439,
    16'd18443,
    16'd18451,
    16'd18457,
    16'd18461,
    16'd18481,
    16'd18493,
    16'd18503,
    16'd18517,
    16'd18521,
    16'd18523,
    16'd18539,
    16'd18541,
    16'd18553,
    16'd18583,
    16'd18587,
    16'd18593,
    16'd18617,
    16'd18637,
    16'd18661,
    16'd18671,
    16'd18679,
    16'd18691,
    16'd18701,
    16'd18713,
    16'd18719,
    16'd18731,
    16'd18743,
    16'd18749,
    16'd18757,
    16'd18773,
    16'd18787,
    16'd18793,
    16'd18797,
    16'd18803,
    16'd18839,
    16'd18859,
    16'd18869,
    16'd18899,
    16'd18911,
    16'd18913,
    16'd18917,
    16'd18919,
    16'd18947,
    16'd18959,
    16'd18973,
    16'd18979,
    16'd19001,
    16'd19009,
    16'd19013,
    16'd19031,
    16'd19037,
    16'd19051,
    16'd19069,
    16'd19073,
    16'd19079,
    16'd19081,
    16'd19087,
    16'd19121,
    16'd19139,
    16'd19141,
    16'd19157,
    16'd19163,
    16'd19181,
    16'd19183,
    16'd19207,
    16'd19211,
    16'd19213,
    16'd19219,
    16'd19231,
    16'd19237,
    16'd19249,
    16'd19259,
    16'd19267,
    16'd19273,
    16'd19289,
    16'd19301,
    16'd19309,
    16'd19319,
    16'd19333,
    16'd19373,
    16'd19379,
    16'd19381,
    16'd19387,
    16'd19391,
    16'd19403,
    16'd19417,
    16'd19421,
    16'd19423,
    16'd19427,
    16'd19429,
    16'd19433,
    16'd19441,
    16'd19447,
    16'd19457,
    16'd19463,
    16'd19469,
    16'd19471,
    16'd19477,
    16'd19483,
    16'd19489,
    16'd19501,
    16'd19507,
    16'd19531,
    16'd19541,
    16'd19543,
    16'd19553,
    16'd19559,
    16'd19571,
    16'd19577,
    16'd19583,
    16'd19597,
    16'd19603,
    16'd19609,
    16'd19661,
    16'd19681,
    16'd19687,
    16'd19697,
    16'd19699,
    16'd19709,
    16'd19717,
    16'd19727,
    16'd19739,
    16'd19751,
    16'd19753,
    16'd19759,
    16'd19763,
    16'd19777,
    16'd19793,
    16'd19801,
    16'd19813,
    16'd19819,
    16'd19841,
    16'd19843,
    16'd19853,
    16'd19861,
    16'd19867,
    16'd19889,
    16'd19891,
    16'd19913,
    16'd19919,
    16'd19927,
    16'd19937,
    16'd19949,
    16'd19961,
    16'd19963,
    16'd19973,
    16'd19979,
    16'd19991,
    16'd19993,
    16'd19997,
    16'd20011,
    16'd20021,
    16'd20023,
    16'd20029,
    16'd20047,
    16'd20051,
    16'd20063,
    16'd20071,
    16'd20089,
    16'd20101,
    16'd20107,
    16'd20113,
    16'd20117,
    16'd20123,
    16'd20129,
    16'd20143,
    16'd20147,
    16'd20149,
    16'd20161,
    16'd20173,
    16'd20177,
    16'd20183,
    16'd20201,
    16'd20219,
    16'd20231,
    16'd20233,
    16'd20249,
    16'd20261,
    16'd20269,
    16'd20287,
    16'd20297,
    16'd20323,
    16'd20327,
    16'd20333,
    16'd20341,
    16'd20347,
    16'd20353,
    16'd20357,
    16'd20359,
    16'd20369,
    16'd20389,
    16'd20393,
    16'd20399,
    16'd20407,
    16'd20411,
    16'd20431,
    16'd20441,
    16'd20443,
    16'd20477,
    16'd20479,
    16'd20483,
    16'd20507,
    16'd20509,
    16'd20521,
    16'd20533,
    16'd20543,
    16'd20549,
    16'd20551,
    16'd20563,
    16'd20593,
    16'd20599,
    16'd20611,
    16'd20627,
    16'd20639,
    16'd20641,
    16'd20663,
    16'd20681,
    16'd20693,
    16'd20707,
    16'd20717,
    16'd20719,
    16'd20731,
    16'd20743,
    16'd20747,
    16'd20749,
    16'd20753,
    16'd20759,
    16'd20771,
    16'd20773,
    16'd20789,
    16'd20807,
    16'd20809,
    16'd20849,
    16'd20857,
    16'd20873,
    16'd20879,
    16'd20887,
    16'd20897,
    16'd20899,
    16'd20903,
    16'd20921,
    16'd20929,
    16'd20939,
    16'd20947,
    16'd20959,
    16'd20963,
    16'd20981,
    16'd20983,
    16'd21001,
    16'd21011,
    16'd21013,
    16'd21017,
    16'd21019,
    16'd21023,
    16'd21031,
    16'd21059,
    16'd21061,
    16'd21067,
    16'd21089,
    16'd21101,
    16'd21107,
    16'd21121,
    16'd21139,
    16'd21143,
    16'd21149,
    16'd21157,
    16'd21163,
    16'd21169,
    16'd21179,
    16'd21187,
    16'd21191,
    16'd21193,
    16'd21211,
    16'd21221,
    16'd21227,
    16'd21247,
    16'd21269,
    16'd21277,
    16'd21283,
    16'd21313,
    16'd21317,
    16'd21319,
    16'd21323,
    16'd21341,
    16'd21347,
    16'd21377,
    16'd21379,
    16'd21383,
    16'd21391,
    16'd21397,
    16'd21401,
    16'd21407,
    16'd21419,
    16'd21433,
    16'd21467,
    16'd21481,
    16'd21487,
    16'd21491,
    16'd21493,
    16'd21499,
    16'd21503,
    16'd21517,
    16'd21521,
    16'd21523,
    16'd21529,
    16'd21557,
    16'd21559,
    16'd21563,
    16'd21569,
    16'd21577,
    16'd21587,
    16'd21589,
    16'd21599,
    16'd21601,
    16'd21611,
    16'd21613,
    16'd21617,
    16'd21647,
    16'd21649,
    16'd21661,
    16'd21673,
    16'd21683,
    16'd21701,
    16'd21713,
    16'd21727,
    16'd21737,
    16'd21739,
    16'd21751,
    16'd21757,
    16'd21767,
    16'd21773,
    16'd21787,
    16'd21799,
    16'd21803,
    16'd21817,
    16'd21821,
    16'd21839,
    16'd21841,
    16'd21851,
    16'd21859,
    16'd21863,
    16'd21871,
    16'd21881,
    16'd21893,
    16'd21911,
    16'd21929,
    16'd21937,
    16'd21943,
    16'd21961,
    16'd21977,
    16'd21991,
    16'd21997,
    16'd22003,
    16'd22013,
    16'd22027,
    16'd22031,
    16'd22037,
    16'd22039,
    16'd22051,
    16'd22063,
    16'd22067,
    16'd22073,
    16'd22079,
    16'd22091,
    16'd22093,
    16'd22109,
    16'd22111,
    16'd22123,
    16'd22129,
    16'd22133,
    16'd22147,
    16'd22153,
    16'd22157,
    16'd22159,
    16'd22171,
    16'd22189,
    16'd22193,
    16'd22229,
    16'd22247,
    16'd22259,
    16'd22271,
    16'd22273,
    16'd22277,
    16'd22279,
    16'd22283,
    16'd22291,
    16'd22303,
    16'd22307,
    16'd22343,
    16'd22349,
    16'd22367,
    16'd22369,
    16'd22381,
    16'd22391,
    16'd22397,
    16'd22409,
    16'd22433,
    16'd22441,
    16'd22447,
    16'd22453,
    16'd22469,
    16'd22481,
    16'd22483,
    16'd22501,
    16'd22511,
    16'd22531,
    16'd22541,
    16'd22543,
    16'd22549,
    16'd22567,
    16'd22571,
    16'd22573,
    16'd22613,
    16'd22619,
    16'd22621,
    16'd22637,
    16'd22639,
    16'd22643,
    16'd22651,
    16'd22669,
    16'd22679,
    16'd22691,
    16'd22697,
    16'd22699,
    16'd22709,
    16'd22717,
    16'd22721,
    16'd22727,
    16'd22739,
    16'd22741,
    16'd22751,
    16'd22769,
    16'd22777,
    16'd22783,
    16'd22787,
    16'd22807,
    16'd22811,
    16'd22817,
    16'd22853,
    16'd22859,
    16'd22861,
    16'd22871,
    16'd22877,
    16'd22901,
    16'd22907,
    16'd22921,
    16'd22937,
    16'd22943,
    16'd22961,
    16'd22963,
    16'd22973,
    16'd22993,
    16'd23003,
    16'd23011,
    16'd23017,
    16'd23021,
    16'd23027,
    16'd23029,
    16'd23039,
    16'd23041,
    16'd23053,
    16'd23057,
    16'd23059,
    16'd23063,
    16'd23071,
    16'd23081,
    16'd23087,
    16'd23099,
    16'd23117,
    16'd23131,
    16'd23143,
    16'd23159,
    16'd23167,
    16'd23173,
    16'd23189,
    16'd23197,
    16'd23201,
    16'd23203,
    16'd23209,
    16'd23227,
    16'd23251,
    16'd23269,
    16'd23279,
    16'd23291,
    16'd23293,
    16'd23297,
    16'd23311,
    16'd23321,
    16'd23327,
    16'd23333,
    16'd23339,
    16'd23357,
    16'd23369,
    16'd23371,
    16'd23399,
    16'd23417,
    16'd23431,
    16'd23447,
    16'd23459,
    16'd23473,
    16'd23497,
    16'd23509,
    16'd23531,
    16'd23537,
    16'd23539,
    16'd23549,
    16'd23557,
    16'd23561,
    16'd23563,
    16'd23567,
    16'd23581,
    16'd23593,
    16'd23599,
    16'd23603,
    16'd23609,
    16'd23623,
    16'd23627,
    16'd23629,
    16'd23633,
    16'd23663,
    16'd23669,
    16'd23671,
    16'd23677,
    16'd23687,
    16'd23689,
    16'd23719,
    16'd23741,
    16'd23743,
    16'd23747,
    16'd23753,
    16'd23761,
    16'd23767,
    16'd23773,
    16'd23789,
    16'd23801,
    16'd23813,
    16'd23819,
    16'd23827,
    16'd23831,
    16'd23833,
    16'd23857,
    16'd23869,
    16'd23873,
    16'd23879,
    16'd23887,
    16'd23893,
    16'd23899,
    16'd23909,
    16'd23911,
    16'd23917,
    16'd23929,
    16'd23957,
    16'd23971,
    16'd23977,
    16'd23981,
    16'd23993,
    16'd24001,
    16'd24007,
    16'd24019,
    16'd24023,
    16'd24029,
    16'd24043,
    16'd24049,
    16'd24061,
    16'd24071,
    16'd24077,
    16'd24083,
    16'd24091,
    16'd24097,
    16'd24103,
    16'd24107,
    16'd24109,
    16'd24113,
    16'd24121,
    16'd24133,
    16'd24137,
    16'd24151,
    16'd24169,
    16'd24179,
    16'd24181,
    16'd24197,
    16'd24203,
    16'd24223,
    16'd24229,
    16'd24239,
    16'd24247,
    16'd24251,
    16'd24281,
    16'd24317,
    16'd24329,
    16'd24337,
    16'd24359,
    16'd24371,
    16'd24373,
    16'd24379,
    16'd24391,
    16'd24407,
    16'd24413,
    16'd24419,
    16'd24421,
    16'd24439,
    16'd24443,
    16'd24469,
    16'd24473,
    16'd24481,
    16'd24499,
    16'd24509,
    16'd24517,
    16'd24527,
    16'd24533,
    16'd24547,
    16'd24551,
    16'd24571,
    16'd24593,
    16'd24611,
    16'd24623,
    16'd24631,
    16'd24659,
    16'd24671,
    16'd24677,
    16'd24683,
    16'd24691,
    16'd24697,
    16'd24709,
    16'd24733,
    16'd24749,
    16'd24763,
    16'd24767,
    16'd24781,
    16'd24793,
    16'd24799,
    16'd24809,
    16'd24821,
    16'd24841,
    16'd24847,
    16'd24851,
    16'd24859,
    16'd24877,
    16'd24889,
    16'd24907,
    16'd24917,
    16'd24919,
    16'd24923,
    16'd24943,
    16'd24953,
    16'd24967,
    16'd24971,
    16'd24977,
    16'd24979,
    16'd24989,
    16'd25013,
    16'd25031,
    16'd25033,
    16'd25037,
    16'd25057,
    16'd25073,
    16'd25087,
    16'd25097,
    16'd25111,
    16'd25117,
    16'd25121,
    16'd25127,
    16'd25147,
    16'd25153,
    16'd25163,
    16'd25169,
    16'd25171,
    16'd25183,
    16'd25189,
    16'd25219,
    16'd25229,
    16'd25237,
    16'd25243,
    16'd25247,
    16'd25253,
    16'd25261,
    16'd25301,
    16'd25303,
    16'd25307,
    16'd25309,
    16'd25321,
    16'd25339,
    16'd25343,
    16'd25349,
    16'd25357,
    16'd25367,
    16'd25373,
    16'd25391,
    16'd25409,
    16'd25411,
    16'd25423,
    16'd25439,
    16'd25447,
    16'd25453,
    16'd25457,
    16'd25463,
    16'd25469,
    16'd25471,
    16'd25523,
    16'd25537,
    16'd25541,
    16'd25561,
    16'd25577,
    16'd25579,
    16'd25583,
    16'd25589,
    16'd25601,
    16'd25603,
    16'd25609,
    16'd25621,
    16'd25633,
    16'd25639,
    16'd25643,
    16'd25657,
    16'd25667,
    16'd25673,
    16'd25679,
    16'd25693,
    16'd25703,
    16'd25717,
    16'd25733,
    16'd25741,
    16'd25747,
    16'd25759,
    16'd25763,
    16'd25771,
    16'd25793,
    16'd25799,
    16'd25801,
    16'd25819,
    16'd25841,
    16'd25847,
    16'd25849,
    16'd25867,
    16'd25873,
    16'd25889,
    16'd25903,
    16'd25913,
    16'd25919,
    16'd25931,
    16'd25933,
    16'd25939,
    16'd25943,
    16'd25951,
    16'd25969,
    16'd25981,
    16'd25997,
    16'd25999,
    16'd26003,
    16'd26017,
    16'd26021,
    16'd26029,
    16'd26041,
    16'd26053,
    16'd26083,
    16'd26099,
    16'd26107,
    16'd26111,
    16'd26113,
    16'd26119,
    16'd26141,
    16'd26153,
    16'd26161,
    16'd26171,
    16'd26177,
    16'd26183,
    16'd26189,
    16'd26203,
    16'd26209,
    16'd26227,
    16'd26237,
    16'd26249,
    16'd26251,
    16'd26261,
    16'd26263,
    16'd26267,
    16'd26293,
    16'd26297,
    16'd26309,
    16'd26317,
    16'd26321,
    16'd26339,
    16'd26347,
    16'd26357,
    16'd26371,
    16'd26387,
    16'd26393,
    16'd26399,
    16'd26407,
    16'd26417,
    16'd26423,
    16'd26431,
    16'd26437,
    16'd26449,
    16'd26459,
    16'd26479,
    16'd26489,
    16'd26497,
    16'd26501,
    16'd26513,
    16'd26539,
    16'd26557,
    16'd26561,
    16'd26573,
    16'd26591,
    16'd26597,
    16'd26627,
    16'd26633,
    16'd26641,
    16'd26647,
    16'd26669,
    16'd26681,
    16'd26683,
    16'd26687,
    16'd26693,
    16'd26699,
    16'd26701,
    16'd26711,
    16'd26713,
    16'd26717,
    16'd26723,
    16'd26729,
    16'd26731,
    16'd26737,
    16'd26759,
    16'd26777,
    16'd26783,
    16'd26801,
    16'd26813,
    16'd26821,
    16'd26833,
    16'd26839,
    16'd26849,
    16'd26861,
    16'd26863,
    16'd26879,
    16'd26881,
    16'd26891,
    16'd26893,
    16'd26903,
    16'd26921,
    16'd26927,
    16'd26947,
    16'd26951,
    16'd26953,
    16'd26959,
    16'd26981,
    16'd26987,
    16'd26993,
    16'd27011,
    16'd27017,
    16'd27031,
    16'd27043,
    16'd27059,
    16'd27061,
    16'd27067,
    16'd27073,
    16'd27077,
    16'd27091,
    16'd27103,
    16'd27107,
    16'd27109,
    16'd27127,
    16'd27143,
    16'd27179,
    16'd27191,
    16'd27197,
    16'd27211,
    16'd27239,
    16'd27241,
    16'd27253,
    16'd27259,
    16'd27271,
    16'd27277,
    16'd27281,
    16'd27283,
    16'd27299,
    16'd27329,
    16'd27337,
    16'd27361,
    16'd27367,
    16'd27397,
    16'd27407,
    16'd27409,
    16'd27427,
    16'd27431,
    16'd27437,
    16'd27449,
    16'd27457,
    16'd27479,
    16'd27481,
    16'd27487,
    16'd27509,
    16'd27527,
    16'd27529,
    16'd27539,
    16'd27541,
    16'd27551,
    16'd27581,
    16'd27583,
    16'd27611,
    16'd27617,
    16'd27631,
    16'd27647,
    16'd27653,
    16'd27673,
    16'd27689,
    16'd27691,
    16'd27697,
    16'd27701,
    16'd27733,
    16'd27737,
    16'd27739,
    16'd27743,
    16'd27749,
    16'd27751,
    16'd27763,
    16'd27767,
    16'd27773,
    16'd27779,
    16'd27791,
    16'd27793,
    16'd27799,
    16'd27803,
    16'd27809,
    16'd27817,
    16'd27823,
    16'd27827,
    16'd27847,
    16'd27851,
    16'd27883,
    16'd27893,
    16'd27901,
    16'd27917,
    16'd27919,
    16'd27941,
    16'd27943,
    16'd27947,
    16'd27953,
    16'd27961,
    16'd27967,
    16'd27983,
    16'd27997,
    16'd28001,
    16'd28019,
    16'd28027,
    16'd28031,
    16'd28051,
    16'd28057,
    16'd28069,
    16'd28081,
    16'd28087,
    16'd28097,
    16'd28099,
    16'd28109,
    16'd28111,
    16'd28123,
    16'd28151,
    16'd28163,
    16'd28181,
    16'd28183,
    16'd28201,
    16'd28211,
    16'd28219,
    16'd28229,
    16'd28277,
    16'd28279,
    16'd28283,
    16'd28289,
    16'd28297,
    16'd28307,
    16'd28309,
    16'd28319,
    16'd28349,
    16'd28351,
    16'd28387,
    16'd28393,
    16'd28403,
    16'd28409,
    16'd28411,
    16'd28429,
    16'd28433,
    16'd28439,
    16'd28447,
    16'd28463,
    16'd28477,
    16'd28493,
    16'd28499,
    16'd28513,
    16'd28517,
    16'd28537,
    16'd28541,
    16'd28547,
    16'd28549,
    16'd28559,
    16'd28571,
    16'd28573,
    16'd28579,
    16'd28591,
    16'd28597,
    16'd28603,
    16'd28607,
    16'd28619,
    16'd28621,
    16'd28627,
    16'd28631,
    16'd28643,
    16'd28649,
    16'd28657,
    16'd28661,
    16'd28663,
    16'd28669,
    16'd28687,
    16'd28697,
    16'd28703,
    16'd28711,
    16'd28723,
    16'd28729,
    16'd28751,
    16'd28753,
    16'd28759,
    16'd28771,
    16'd28789,
    16'd28793,
    16'd28807,
    16'd28813,
    16'd28817,
    16'd28837,
    16'd28843,
    16'd28859,
    16'd28867,
    16'd28871,
    16'd28879,
    16'd28901,
    16'd28909,
    16'd28921,
    16'd28927,
    16'd28933,
    16'd28949,
    16'd28961,
    16'd28979,
    16'd29009,
    16'd29017,
    16'd29021,
    16'd29023,
    16'd29027,
    16'd29033,
    16'd29059,
    16'd29063,
    16'd29077,
    16'd29101,
    16'd29123,
    16'd29129,
    16'd29131,
    16'd29137,
    16'd29147,
    16'd29153,
    16'd29167,
    16'd29173,
    16'd29179,
    16'd29191,
    16'd29201,
    16'd29207,
    16'd29209,
    16'd29221,
    16'd29231,
    16'd29243,
    16'd29251,
    16'd29269,
    16'd29287,
    16'd29297,
    16'd29303,
    16'd29311,
    16'd29327,
    16'd29333,
    16'd29339,
    16'd29347,
    16'd29363,
    16'd29383,
    16'd29387,
    16'd29389,
    16'd29399,
    16'd29401,
    16'd29411,
    16'd29423,
    16'd29429,
    16'd29437,
    16'd29443,
    16'd29453,
    16'd29473,
    16'd29483,
    16'd29501,
    16'd29527,
    16'd29531,
    16'd29537,
    16'd29567,
    16'd29569,
    16'd29573,
    16'd29581,
    16'd29587,
    16'd29599,
    16'd29611,
    16'd29629,
    16'd29633,
    16'd29641,
    16'd29663,
    16'd29669,
    16'd29671,
    16'd29683,
    16'd29717,
    16'd29723,
    16'd29741,
    16'd29753,
    16'd29759,
    16'd29761,
    16'd29789,
    16'd29803,
    16'd29819,
    16'd29833,
    16'd29837,
    16'd29851,
    16'd29863,
    16'd29867,
    16'd29873,
    16'd29879,
    16'd29881,
    16'd29917,
    16'd29921,
    16'd29927,
    16'd29947,
    16'd29959,
    16'd29983,
    16'd29989,
    16'd30011,
    16'd30013,
    16'd30029,
    16'd30047,
    16'd30059,
    16'd30071,
    16'd30089,
    16'd30091,
    16'd30097,
    16'd30103,
    16'd30109,
    16'd30113,
    16'd30119,
    16'd30133,
    16'd30137,
    16'd30139,
    16'd30161,
    16'd30169,
    16'd30181,
    16'd30187,
    16'd30197,
    16'd30203,
    16'd30211,
    16'd30223,
    16'd30241,
    16'd30253,
    16'd30259,
    16'd30269,
    16'd30271,
    16'd30293,
    16'd30307,
    16'd30313,
    16'd30319,
    16'd30323,
    16'd30341,
    16'd30347,
    16'd30367,
    16'd30389,
    16'd30391,
    16'd30403,
    16'd30427,
    16'd30431,
    16'd30449,
    16'd30467,
    16'd30469,
    16'd30491,
    16'd30493,
    16'd30497,
    16'd30509,
    16'd30517,
    16'd30529,
    16'd30539,
    16'd30553,
    16'd30557,
    16'd30559,
    16'd30577,
    16'd30593,
    16'd30631,
    16'd30637,
    16'd30643,
    16'd30649,
    16'd30661,
    16'd30671,
    16'd30677,
    16'd30689,
    16'd30697,
    16'd30703,
    16'd30707,
    16'd30713,
    16'd30727,
    16'd30757,
    16'd30763,
    16'd30773,
    16'd30781,
    16'd30803,
    16'd30809,
    16'd30817,
    16'd30829,
    16'd30839,
    16'd30841,
    16'd30851,
    16'd30853,
    16'd30859,
    16'd30869,
    16'd30871,
    16'd30881,
    16'd30893,
    16'd30911,
    16'd30931,
    16'd30937,
    16'd30941,
    16'd30949,
    16'd30971,
    16'd30977,
    16'd30983,
    16'd31013,
    16'd31019,
    16'd31033,
    16'd31039,
    16'd31051,
    16'd31063,
    16'd31069,
    16'd31079,
    16'd31081,
    16'd31091,
    16'd31121,
    16'd31123,
    16'd31139,
    16'd31147,
    16'd31151,
    16'd31153,
    16'd31159,
    16'd31177,
    16'd31181,
    16'd31183,
    16'd31189,
    16'd31193,
    16'd31219,
    16'd31223,
    16'd31231,
    16'd31237,
    16'd31247,
    16'd31249,
    16'd31253,
    16'd31259,
    16'd31267,
    16'd31271,
    16'd31277,
    16'd31307,
    16'd31319,
    16'd31321,
    16'd31327,
    16'd31333,
    16'd31337,
    16'd31357,
    16'd31379,
    16'd31387,
    16'd31391,
    16'd31393,
    16'd31397,
    16'd31469,
    16'd31477,
    16'd31481,
    16'd31489,
    16'd31511,
    16'd31513,
    16'd31517,
    16'd31531,
    16'd31541,
    16'd31543,
    16'd31547,
    16'd31567,
    16'd31573,
    16'd31583,
    16'd31601,
    16'd31607,
    16'd31627,
    16'd31643,
    16'd31649,
    16'd31657,
    16'd31663,
    16'd31667,
    16'd31687,
    16'd31699,
    16'd31721,
    16'd31723,
    16'd31727,
    16'd31729,
    16'd31741,
    16'd31751,
    16'd31769,
    16'd31771,
    16'd31793,
    16'd31799,
    16'd31817,
    16'd31847,
    16'd31849,
    16'd31859,
    16'd31873,
    16'd31883,
    16'd31891,
    16'd31907,
    16'd31957,
    16'd31963,
    16'd31973,
    16'd31981,
    16'd31991,
    16'd32003,
    16'd32009,
    16'd32027,
    16'd32029,
    16'd32051,
    16'd32057,
    16'd32059,
    16'd32063,
    16'd32069,
    16'd32077,
    16'd32083,
    16'd32089,
    16'd32099,
    16'd32117,
    16'd32119,
    16'd32141,
    16'd32143,
    16'd32159,
    16'd32173,
    16'd32183,
    16'd32189,
    16'd32191,
    16'd32203,
    16'd32213,
    16'd32233,
    16'd32237,
    16'd32251,
    16'd32257,
    16'd32261,
    16'd32297,
    16'd32299,
    16'd32303,
    16'd32309,
    16'd32321,
    16'd32323,
    16'd32327,
    16'd32341,
    16'd32353,
    16'd32359,
    16'd32363,
    16'd32369,
    16'd32371,
    16'd32377,
    16'd32381,
    16'd32401,
    16'd32411,
    16'd32413,
    16'd32423,
    16'd32429,
    16'd32441,
    16'd32443,
    16'd32467,
    16'd32479,
    16'd32491,
    16'd32497,
    16'd32503,
    16'd32507,
    16'd32531,
    16'd32533,
    16'd32537,
    16'd32561,
    16'd32563,
    16'd32569,
    16'd32573,
    16'd32579,
    16'd32587,
    16'd32603,
    16'd32609,
    16'd32611,
    16'd32621,
    16'd32633,
    16'd32647,
    16'd32653,
    16'd32687,
    16'd32693,
    16'd32707,
    16'd32713,
    16'd32717,
    16'd32719,
    16'd32749,
    16'd32771,
    16'd32779,
    16'd32783,
    16'd32789,
    16'd32797,
    16'd32801,
    16'd32803,
    16'd32831,
    16'd32833,
    16'd32839,
    16'd32843,
    16'd32869,
    16'd32887,
    16'd32909,
    16'd32911,
    16'd32917,
    16'd32933,
    16'd32939,
    16'd32941,
    16'd32957,
    16'd32969,
    16'd32971,
    16'd32983,
    16'd32987,
    16'd32993,
    16'd32999,
    16'd33013,
    16'd33023,
    16'd33029,
    16'd33037,
    16'd33049,
    16'd33053,
    16'd33071,
    16'd33073,
    16'd33083,
    16'd33091,
    16'd33107,
    16'd33113,
    16'd33119,
    16'd33149,
    16'd33151,
    16'd33161,
    16'd33179,
    16'd33181,
    16'd33191,
    16'd33199,
    16'd33203,
    16'd33211,
    16'd33223,
    16'd33247,
    16'd33287,
    16'd33289,
    16'd33301,
    16'd33311,
    16'd33317,
    16'd33329,
    16'd33331,
    16'd33343,
    16'd33347,
    16'd33349,
    16'd33353,
    16'd33359,
    16'd33377,
    16'd33391,
    16'd33403,
    16'd33409,
    16'd33413,
    16'd33427,
    16'd33457,
    16'd33461,
    16'd33469,
    16'd33479,
    16'd33487,
    16'd33493,
    16'd33503,
    16'd33521,
    16'd33529,
    16'd33533,
    16'd33547,
    16'd33563,
    16'd33569,
    16'd33577,
    16'd33581,
    16'd33587,
    16'd33589,
    16'd33599,
    16'd33601,
    16'd33613,
    16'd33617,
    16'd33619,
    16'd33623,
    16'd33629,
    16'd33637,
    16'd33641,
    16'd33647,
    16'd33679,
    16'd33703,
    16'd33713,
    16'd33721,
    16'd33739,
    16'd33749,
    16'd33751,
    16'd33757,
    16'd33767,
    16'd33769,
    16'd33773,
    16'd33791,
    16'd33797,
    16'd33809,
    16'd33811,
    16'd33827,
    16'd33829,
    16'd33851,
    16'd33857,
    16'd33863,
    16'd33871,
    16'd33889,
    16'd33893,
    16'd33911,
    16'd33923,
    16'd33931,
    16'd33937,
    16'd33941,
    16'd33961,
    16'd33967,
    16'd33997,
    16'd34019,
    16'd34031,
    16'd34033,
    16'd34039,
    16'd34057,
    16'd34061,
    16'd34123,
    16'd34127,
    16'd34129,
    16'd34141,
    16'd34147,
    16'd34157,
    16'd34159,
    16'd34171,
    16'd34183,
    16'd34211,
    16'd34213,
    16'd34217,
    16'd34231,
    16'd34253,
    16'd34259,
    16'd34261,
    16'd34267,
    16'd34273,
    16'd34283,
    16'd34297,
    16'd34301,
    16'd34303,
    16'd34313,
    16'd34319,
    16'd34327,
    16'd34337,
    16'd34351,
    16'd34361,
    16'd34367,
    16'd34369,
    16'd34381,
    16'd34403,
    16'd34421,
    16'd34429,
    16'd34439,
    16'd34457,
    16'd34469,
    16'd34471,
    16'd34483,
    16'd34487,
    16'd34499,
    16'd34501,
    16'd34511,
    16'd34513,
    16'd34519,
    16'd34537,
    16'd34543,
    16'd34549,
    16'd34583,
    16'd34589,
    16'd34591,
    16'd34603,
    16'd34607,
    16'd34613,
    16'd34631,
    16'd34649,
    16'd34651,
    16'd34667,
    16'd34673,
    16'd34679,
    16'd34687,
    16'd34693,
    16'd34703,
    16'd34721,
    16'd34729,
    16'd34739,
    16'd34747,
    16'd34757,
    16'd34759,
    16'd34763,
    16'd34781,
    16'd34807,
    16'd34819,
    16'd34841,
    16'd34843,
    16'd34847,
    16'd34849,
    16'd34871,
    16'd34877,
    16'd34883,
    16'd34897,
    16'd34913,
    16'd34919,
    16'd34939,
    16'd34949,
    16'd34961,
    16'd34963,
    16'd34981,
    16'd35023,
    16'd35027,
    16'd35051,
    16'd35053,
    16'd35059,
    16'd35069,
    16'd35081,
    16'd35083,
    16'd35089,
    16'd35099,
    16'd35107,
    16'd35111,
    16'd35117,
    16'd35129,
    16'd35141,
    16'd35149,
    16'd35153,
    16'd35159,
    16'd35171,
    16'd35201,
    16'd35221,
    16'd35227,
    16'd35251,
    16'd35257,
    16'd35267,
    16'd35279,
    16'd35281,
    16'd35291,
    16'd35311,
    16'd35317,
    16'd35323,
    16'd35327,
    16'd35339,
    16'd35353,
    16'd35363,
    16'd35381,
    16'd35393,
    16'd35401,
    16'd35407,
    16'd35419,
    16'd35423,
    16'd35437,
    16'd35447,
    16'd35449,
    16'd35461,
    16'd35491,
    16'd35507,
    16'd35509,
    16'd35521,
    16'd35527,
    16'd35531,
    16'd35533,
    16'd35537,
    16'd35543,
    16'd35569,
    16'd35573,
    16'd35591,
    16'd35593,
    16'd35597,
    16'd35603,
    16'd35617,
    16'd35671,
    16'd35677,
    16'd35729,
    16'd35731,
    16'd35747,
    16'd35753,
    16'd35759,
    16'd35771,
    16'd35797,
    16'd35801,
    16'd35803,
    16'd35809,
    16'd35831,
    16'd35837,
    16'd35839,
    16'd35851,
    16'd35863,
    16'd35869,
    16'd35879,
    16'd35897,
    16'd35899,
    16'd35911,
    16'd35923,
    16'd35933,
    16'd35951,
    16'd35963,
    16'd35969,
    16'd35977,
    16'd35983,
    16'd35993,
    16'd35999,
    16'd36007,
    16'd36011,
    16'd36013,
    16'd36017,
    16'd36037,
    16'd36061,
    16'd36067,
    16'd36073,
    16'd36083,
    16'd36097,
    16'd36107,
    16'd36109,
    16'd36131,
    16'd36137,
    16'd36151,
    16'd36161,
    16'd36187,
    16'd36191,
    16'd36209,
    16'd36217,
    16'd36229,
    16'd36241,
    16'd36251,
    16'd36263,
    16'd36269,
    16'd36277,
    16'd36293,
    16'd36299,
    16'd36307,
    16'd36313,
    16'd36319,
    16'd36341,
    16'd36343,
    16'd36353,
    16'd36373,
    16'd36383,
    16'd36389,
    16'd36433,
    16'd36451,
    16'd36457,
    16'd36467,
    16'd36469,
    16'd36473,
    16'd36479,
    16'd36493,
    16'd36497,
    16'd36523,
    16'd36527,
    16'd36529,
    16'd36541,
    16'd36551,
    16'd36559,
    16'd36563,
    16'd36571,
    16'd36583,
    16'd36587,
    16'd36599,
    16'd36607,
    16'd36629,
    16'd36637,
    16'd36643,
    16'd36653,
    16'd36671,
    16'd36677,
    16'd36683,
    16'd36691,
    16'd36697,
    16'd36709,
    16'd36713,
    16'd36721,
    16'd36739,
    16'd36749,
    16'd36761,
    16'd36767,
    16'd36779,
    16'd36781,
    16'd36787,
    16'd36791,
    16'd36793,
    16'd36809,
    16'd36821,
    16'd36833,
    16'd36847,
    16'd36857,
    16'd36871,
    16'd36877,
    16'd36887,
    16'd36899,
    16'd36901,
    16'd36913,
    16'd36919,
    16'd36923,
    16'd36929,
    16'd36931,
    16'd36943,
    16'd36947,
    16'd36973,
    16'd36979,
    16'd36997,
    16'd37003,
    16'd37013,
    16'd37019,
    16'd37021,
    16'd37039,
    16'd37049,
    16'd37057,
    16'd37061,
    16'd37087,
    16'd37097,
    16'd37117,
    16'd37123,
    16'd37139,
    16'd37159,
    16'd37171,
    16'd37181,
    16'd37189,
    16'd37199,
    16'd37201,
    16'd37217,
    16'd37223,
    16'd37243,
    16'd37253,
    16'd37273,
    16'd37277,
    16'd37307,
    16'd37309,
    16'd37313,
    16'd37321,
    16'd37337,
    16'd37339,
    16'd37357,
    16'd37361,
    16'd37363,
    16'd37369,
    16'd37379,
    16'd37397,
    16'd37409,
    16'd37423,
    16'd37441,
    16'd37447,
    16'd37463,
    16'd37483,
    16'd37489,
    16'd37493,
    16'd37501,
    16'd37507,
    16'd37511,
    16'd37517,
    16'd37529,
    16'd37537,
    16'd37547,
    16'd37549,
    16'd37561,
    16'd37567,
    16'd37571,
    16'd37573,
    16'd37579,
    16'd37589,
    16'd37591,
    16'd37607,
    16'd37619,
    16'd37633,
    16'd37643,
    16'd37649,
    16'd37657,
    16'd37663,
    16'd37691,
    16'd37693,
    16'd37699,
    16'd37717,
    16'd37747,
    16'd37781,
    16'd37783,
    16'd37799,
    16'd37811,
    16'd37813,
    16'd37831,
    16'd37847,
    16'd37853,
    16'd37861,
    16'd37871,
    16'd37879,
    16'd37889,
    16'd37897,
    16'd37907,
    16'd37951,
    16'd37957,
    16'd37963,
    16'd37967,
    16'd37987,
    16'd37991,
    16'd37993,
    16'd37997,
    16'd38011,
    16'd38039,
    16'd38047,
    16'd38053,
    16'd38069,
    16'd38083,
    16'd38113,
    16'd38119,
    16'd38149,
    16'd38153,
    16'd38167,
    16'd38177,
    16'd38183,
    16'd38189,
    16'd38197,
    16'd38201,
    16'd38219,
    16'd38231,
    16'd38237,
    16'd38239,
    16'd38261,
    16'd38273,
    16'd38281,
    16'd38287,
    16'd38299,
    16'd38303,
    16'd38317,
    16'd38321,
    16'd38327,
    16'd38329,
    16'd38333,
    16'd38351,
    16'd38371,
    16'd38377,
    16'd38393,
    16'd38431,
    16'd38447,
    16'd38449,
    16'd38453,
    16'd38459,
    16'd38461,
    16'd38501,
    16'd38543,
    16'd38557,
    16'd38561,
    16'd38567,
    16'd38569,
    16'd38593,
    16'd38603,
    16'd38609,
    16'd38611,
    16'd38629,
    16'd38639,
    16'd38651,
    16'd38653,
    16'd38669,
    16'd38671,
    16'd38677,
    16'd38693,
    16'd38699,
    16'd38707,
    16'd38711,
    16'd38713,
    16'd38723,
    16'd38729,
    16'd38737,
    16'd38747,
    16'd38749,
    16'd38767,
    16'd38783,
    16'd38791,
    16'd38803,
    16'd38821,
    16'd38833,
    16'd38839,
    16'd38851,
    16'd38861,
    16'd38867,
    16'd38873,
    16'd38891,
    16'd38903,
    16'd38917,
    16'd38921,
    16'd38923,
    16'd38933,
    16'd38953,
    16'd38959,
    16'd38971,
    16'd38977,
    16'd38993,
    16'd39019,
    16'd39023,
    16'd39041,
    16'd39043,
    16'd39047,
    16'd39079,
    16'd39089,
    16'd39097,
    16'd39103,
    16'd39107,
    16'd39113,
    16'd39119,
    16'd39133,
    16'd39139,
    16'd39157,
    16'd39161,
    16'd39163,
    16'd39181,
    16'd39191,
    16'd39199,
    16'd39209,
    16'd39217,
    16'd39227,
    16'd39229,
    16'd39233,
    16'd39239,
    16'd39241,
    16'd39251,
    16'd39293,
    16'd39301,
    16'd39313,
    16'd39317,
    16'd39323,
    16'd39341,
    16'd39343,
    16'd39359,
    16'd39367,
    16'd39371,
    16'd39373,
    16'd39383,
    16'd39397,
    16'd39409,
    16'd39419,
    16'd39439,
    16'd39443,
    16'd39451,
    16'd39461,
    16'd39499,
    16'd39503,
    16'd39509,
    16'd39511,
    16'd39521,
    16'd39541,
    16'd39551,
    16'd39563,
    16'd39569,
    16'd39581,
    16'd39607,
    16'd39619,
    16'd39623,
    16'd39631,
    16'd39659,
    16'd39667,
    16'd39671,
    16'd39679,
    16'd39703,
    16'd39709,
    16'd39719,
    16'd39727,
    16'd39733,
    16'd39749,
    16'd39761,
    16'd39769,
    16'd39779,
    16'd39791,
    16'd39799,
    16'd39821,
    16'd39827,
    16'd39829,
    16'd39839,
    16'd39841,
    16'd39847,
    16'd39857,
    16'd39863,
    16'd39869,
    16'd39877,
    16'd39883,
    16'd39887,
    16'd39901,
    16'd39929,
    16'd39937,
    16'd39953,
    16'd39971,
    16'd39979,
    16'd39983,
    16'd39989,
    16'd40009,
    16'd40013,
    16'd40031,
    16'd40037,
    16'd40039,
    16'd40063,
    16'd40087,
    16'd40093,
    16'd40099,
    16'd40111,
    16'd40123,
    16'd40127,
    16'd40129,
    16'd40151,
    16'd40153,
    16'd40163,
    16'd40169,
    16'd40177,
    16'd40189,
    16'd40193,
    16'd40213,
    16'd40231,
    16'd40237,
    16'd40241,
    16'd40253,
    16'd40277,
    16'd40283,
    16'd40289,
    16'd40343,
    16'd40351,
    16'd40357,
    16'd40361,
    16'd40387,
    16'd40423,
    16'd40427,
    16'd40429,
    16'd40433,
    16'd40459,
    16'd40471,
    16'd40483,
    16'd40487,
    16'd40493,
    16'd40499,
    16'd40507,
    16'd40519,
    16'd40529,
    16'd40531,
    16'd40543,
    16'd40559,
    16'd40577,
    16'd40583,
    16'd40591,
    16'd40597,
    16'd40609,
    16'd40627,
    16'd40637,
    16'd40639,
    16'd40693,
    16'd40697,
    16'd40699,
    16'd40709,
    16'd40739,
    16'd40751,
    16'd40759,
    16'd40763,
    16'd40771,
    16'd40787,
    16'd40801,
    16'd40813,
    16'd40819,
    16'd40823,
    16'd40829,
    16'd40841,
    16'd40847,
    16'd40849,
    16'd40853,
    16'd40867,
    16'd40879,
    16'd40883,
    16'd40897,
    16'd40903,
    16'd40927,
    16'd40933,
    16'd40939,
    16'd40949,
    16'd40961,
    16'd40973,
    16'd40993,
    16'd41011,
    16'd41017,
    16'd41023,
    16'd41039,
    16'd41047,
    16'd41051,
    16'd41057,
    16'd41077,
    16'd41081,
    16'd41113,
    16'd41117,
    16'd41131,
    16'd41141,
    16'd41143,
    16'd41149,
    16'd41161,
    16'd41177,
    16'd41179,
    16'd41183,
    16'd41189,
    16'd41201,
    16'd41203,
    16'd41213,
    16'd41221,
    16'd41227,
    16'd41231,
    16'd41233,
    16'd41243,
    16'd41257,
    16'd41263,
    16'd41269,
    16'd41281,
    16'd41299,
    16'd41333,
    16'd41341,
    16'd41351,
    16'd41357,
    16'd41381,
    16'd41387,
    16'd41389,
    16'd41399,
    16'd41411,
    16'd41413,
    16'd41443,
    16'd41453,
    16'd41467,
    16'd41479,
    16'd41491,
    16'd41507,
    16'd41513,
    16'd41519,
    16'd41521,
    16'd41539,
    16'd41543,
    16'd41549,
    16'd41579,
    16'd41593,
    16'd41597,
    16'd41603,
    16'd41609,
    16'd41611,
    16'd41617,
    16'd41621,
    16'd41627,
    16'd41641,
    16'd41647,
    16'd41651,
    16'd41659,
    16'd41669,
    16'd41681,
    16'd41687,
    16'd41719,
    16'd41729,
    16'd41737,
    16'd41759,
    16'd41761,
    16'd41771,
    16'd41777,
    16'd41801,
    16'd41809,
    16'd41813,
    16'd41843,
    16'd41849,
    16'd41851,
    16'd41863,
    16'd41879,
    16'd41887,
    16'd41893,
    16'd41897,
    16'd41903,
    16'd41911,
    16'd41927,
    16'd41941,
    16'd41947,
    16'd41953,
    16'd41957,
    16'd41959,
    16'd41969,
    16'd41981,
    16'd41983,
    16'd41999,
    16'd42013,
    16'd42017,
    16'd42019,
    16'd42023,
    16'd42043,
    16'd42061,
    16'd42071,
    16'd42073,
    16'd42083,
    16'd42089,
    16'd42101,
    16'd42131,
    16'd42139,
    16'd42157,
    16'd42169,
    16'd42179,
    16'd42181,
    16'd42187,
    16'd42193,
    16'd42197,
    16'd42209,
    16'd42221,
    16'd42223,
    16'd42227,
    16'd42239,
    16'd42257,
    16'd42281,
    16'd42283,
    16'd42293,
    16'd42299,
    16'd42307,
    16'd42323,
    16'd42331,
    16'd42337,
    16'd42349,
    16'd42359,
    16'd42373,
    16'd42379,
    16'd42391,
    16'd42397,
    16'd42403,
    16'd42407,
    16'd42409,
    16'd42433,
    16'd42437,
    16'd42443,
    16'd42451,
    16'd42457,
    16'd42461,
    16'd42463,
    16'd42467,
    16'd42473,
    16'd42487,
    16'd42491,
    16'd42499,
    16'd42509,
    16'd42533,
    16'd42557,
    16'd42569,
    16'd42571,
    16'd42577,
    16'd42589,
    16'd42611,
    16'd42641,
    16'd42643,
    16'd42649,
    16'd42667,
    16'd42677,
    16'd42683,
    16'd42689,
    16'd42697,
    16'd42701,
    16'd42703,
    16'd42709,
    16'd42719,
    16'd42727,
    16'd42737,
    16'd42743,
    16'd42751,
    16'd42767,
    16'd42773,
    16'd42787,
    16'd42793,
    16'd42797,
    16'd42821,
    16'd42829,
    16'd42839,
    16'd42841,
    16'd42853,
    16'd42859,
    16'd42863,
    16'd42899,
    16'd42901,
    16'd42923,
    16'd42929,
    16'd42937,
    16'd42943,
    16'd42953,
    16'd42961,
    16'd42967,
    16'd42979,
    16'd42989,
    16'd43003,
    16'd43013,
    16'd43019,
    16'd43037,
    16'd43049,
    16'd43051,
    16'd43063,
    16'd43067,
    16'd43093,
    16'd43103,
    16'd43117,
    16'd43133,
    16'd43151,
    16'd43159,
    16'd43177,
    16'd43189,
    16'd43201,
    16'd43207,
    16'd43223,
    16'd43237,
    16'd43261,
    16'd43271,
    16'd43283,
    16'd43291,
    16'd43313,
    16'd43319,
    16'd43321,
    16'd43331,
    16'd43391,
    16'd43397,
    16'd43399,
    16'd43403,
    16'd43411,
    16'd43427,
    16'd43441,
    16'd43451,
    16'd43457,
    16'd43481,
    16'd43487,
    16'd43499,
    16'd43517,
    16'd43541,
    16'd43543,
    16'd43573,
    16'd43577,
    16'd43579,
    16'd43591,
    16'd43597,
    16'd43607,
    16'd43609,
    16'd43613,
    16'd43627,
    16'd43633,
    16'd43649,
    16'd43651,
    16'd43661,
    16'd43669,
    16'd43691,
    16'd43711,
    16'd43717,
    16'd43721,
    16'd43753,
    16'd43759,
    16'd43777,
    16'd43781,
    16'd43783,
    16'd43787,
    16'd43789,
    16'd43793,
    16'd43801,
    16'd43853,
    16'd43867,
    16'd43889,
    16'd43891,
    16'd43913,
    16'd43933,
    16'd43943,
    16'd43951,
    16'd43961,
    16'd43963,
    16'd43969,
    16'd43973,
    16'd43987,
    16'd43991,
    16'd43997,
    16'd44017,
    16'd44021,
    16'd44027,
    16'd44029,
    16'd44041,
    16'd44053,
    16'd44059,
    16'd44071,
    16'd44087,
    16'd44089,
    16'd44101,
    16'd44111,
    16'd44119,
    16'd44123,
    16'd44129,
    16'd44131,
    16'd44159,
    16'd44171,
    16'd44179,
    16'd44189,
    16'd44201,
    16'd44203,
    16'd44207,
    16'd44221,
    16'd44249,
    16'd44257,
    16'd44263,
    16'd44267,
    16'd44269,
    16'd44273,
    16'd44279,
    16'd44281,
    16'd44293,
    16'd44351,
    16'd44357,
    16'd44371,
    16'd44381,
    16'd44383,
    16'd44389,
    16'd44417,
    16'd44449,
    16'd44453,
    16'd44483,
    16'd44491,
    16'd44497,
    16'd44501,
    16'd44507,
    16'd44519,
    16'd44531,
    16'd44533,
    16'd44537,
    16'd44543,
    16'd44549,
    16'd44563,
    16'd44579,
    16'd44587,
    16'd44617,
    16'd44621,
    16'd44623,
    16'd44633,
    16'd44641,
    16'd44647,
    16'd44651,
    16'd44657,
    16'd44683,
    16'd44687,
    16'd44699,
    16'd44701,
    16'd44711,
    16'd44729,
    16'd44741,
    16'd44753,
    16'd44771,
    16'd44773,
    16'd44777,
    16'd44789,
    16'd44797,
    16'd44809,
    16'd44819,
    16'd44839,
    16'd44843,
    16'd44851,
    16'd44867,
    16'd44879,
    16'd44887,
    16'd44893,
    16'd44909,
    16'd44917,
    16'd44927,
    16'd44939,
    16'd44953,
    16'd44959,
    16'd44963,
    16'd44971,
    16'd44983,
    16'd44987,
    16'd45007,
    16'd45013,
    16'd45053,
    16'd45061,
    16'd45077,
    16'd45083,
    16'd45119,
    16'd45121,
    16'd45127,
    16'd45131,
    16'd45137,
    16'd45139,
    16'd45161,
    16'd45179,
    16'd45181,
    16'd45191,
    16'd45197,
    16'd45233,
    16'd45247,
    16'd45259,
    16'd45263,
    16'd45281,
    16'd45289,
    16'd45293,
    16'd45307,
    16'd45317,
    16'd45319,
    16'd45329,
    16'd45337,
    16'd45341,
    16'd45343,
    16'd45361,
    16'd45377,
    16'd45389,
    16'd45403,
    16'd45413,
    16'd45427,
    16'd45433,
    16'd45439,
    16'd45481,
    16'd45491,
    16'd45497,
    16'd45503,
    16'd45523,
    16'd45533,
    16'd45541,
    16'd45553,
    16'd45557,
    16'd45569,
    16'd45587,
    16'd45589,
    16'd45599,
    16'd45613,
    16'd45631,
    16'd45641,
    16'd45659,
    16'd45667,
    16'd45673,
    16'd45677,
    16'd45691,
    16'd45697,
    16'd45707,
    16'd45737,
    16'd45751,
    16'd45757,
    16'd45763,
    16'd45767,
    16'd45779,
    16'd45817,
    16'd45821,
    16'd45823,
    16'd45827,
    16'd45833,
    16'd45841,
    16'd45853,
    16'd45863,
    16'd45869,
    16'd45887,
    16'd45893,
    16'd45943,
    16'd45949,
    16'd45953,
    16'd45959,
    16'd45971,
    16'd45979,
    16'd45989,
    16'd46021,
    16'd46027,
    16'd46049,
    16'd46051,
    16'd46061,
    16'd46073,
    16'd46091,
    16'd46093,
    16'd46099,
    16'd46103,
    16'd46133,
    16'd46141,
    16'd46147,
    16'd46153,
    16'd46171,
    16'd46181,
    16'd46183,
    16'd46187,
    16'd46199,
    16'd46219,
    16'd46229,
    16'd46237,
    16'd46261,
    16'd46271,
    16'd46273,
    16'd46279,
    16'd46301,
    16'd46307,
    16'd46309,
    16'd46327,
    16'd46337,
    16'd46349,
    16'd46351,
    16'd46381,
    16'd46399,
    16'd46411,
    16'd46439,
    16'd46441,
    16'd46447,
    16'd46451,
    16'd46457,
    16'd46471,
    16'd46477,
    16'd46489,
    16'd46499,
    16'd46507,
    16'd46511,
    16'd46523,
    16'd46549,
    16'd46559,
    16'd46567,
    16'd46573,
    16'd46589,
    16'd46591,
    16'd46601,
    16'd46619,
    16'd46633,
    16'd46639,
    16'd46643,
    16'd46649,
    16'd46663,
    16'd46679,
    16'd46681,
    16'd46687,
    16'd46691,
    16'd46703,
    16'd46723,
    16'd46727,
    16'd46747,
    16'd46751,
    16'd46757,
    16'd46769,
    16'd46771,
    16'd46807,
    16'd46811,
    16'd46817,
    16'd46819,
    16'd46829,
    16'd46831,
    16'd46853,
    16'd46861,
    16'd46867,
    16'd46877,
    16'd46889,
    16'd46901,
    16'd46919,
    16'd46933,
    16'd46957,
    16'd46993,
    16'd46997,
    16'd47017,
    16'd47041,
    16'd47051,
    16'd47057,
    16'd47059,
    16'd47087,
    16'd47093,
    16'd47111,
    16'd47119,
    16'd47123,
    16'd47129,
    16'd47137,
    16'd47143,
    16'd47147,
    16'd47149,
    16'd47161,
    16'd47189,
    16'd47207,
    16'd47221,
    16'd47237,
    16'd47251,
    16'd47269,
    16'd47279,
    16'd47287,
    16'd47293,
    16'd47297,
    16'd47303,
    16'd47309,
    16'd47317,
    16'd47339,
    16'd47351,
    16'd47353,
    16'd47363,
    16'd47381,
    16'd47387,
    16'd47389,
    16'd47407,
    16'd47417,
    16'd47419,
    16'd47431,
    16'd47441,
    16'd47459,
    16'd47491,
    16'd47497,
    16'd47501,
    16'd47507,
    16'd47513,
    16'd47521,
    16'd47527,
    16'd47533,
    16'd47543,
    16'd47563,
    16'd47569,
    16'd47581,
    16'd47591,
    16'd47599,
    16'd47609,
    16'd47623,
    16'd47629,
    16'd47639,
    16'd47653,
    16'd47657,
    16'd47659,
    16'd47681,
    16'd47699,
    16'd47701,
    16'd47711,
    16'd47713,
    16'd47717,
    16'd47737,
    16'd47741,
    16'd47743,
    16'd47777,
    16'd47779,
    16'd47791,
    16'd47797,
    16'd47807,
    16'd47809,
    16'd47819,
    16'd47837,
    16'd47843,
    16'd47857,
    16'd47869,
    16'd47881,
    16'd47903,
    16'd47911,
    16'd47917,
    16'd47933,
    16'd47939,
    16'd47947,
    16'd47951,
    16'd47963,
    16'd47969,
    16'd47977,
    16'd47981,
    16'd48017,
    16'd48023,
    16'd48029,
    16'd48049,
    16'd48073,
    16'd48079,
    16'd48091,
    16'd48109,
    16'd48119,
    16'd48121,
    16'd48131,
    16'd48157,
    16'd48163,
    16'd48179,
    16'd48187,
    16'd48193,
    16'd48197,
    16'd48221,
    16'd48239,
    16'd48247,
    16'd48259,
    16'd48271,
    16'd48281,
    16'd48299,
    16'd48311,
    16'd48313,
    16'd48337,
    16'd48341,
    16'd48353,
    16'd48371,
    16'd48383,
    16'd48397,
    16'd48407,
    16'd48409,
    16'd48413,
    16'd48437,
    16'd48449,
    16'd48463,
    16'd48473,
    16'd48479,
    16'd48481,
    16'd48487,
    16'd48491,
    16'd48497,
    16'd48523,
    16'd48527,
    16'd48533,
    16'd48539,
    16'd48541,
    16'd48563,
    16'd48571,
    16'd48589,
    16'd48593,
    16'd48611,
    16'd48619,
    16'd48623,
    16'd48647,
    16'd48649,
    16'd48661,
    16'd48673,
    16'd48677,
    16'd48679,
    16'd48731,
    16'd48733,
    16'd48751,
    16'd48757,
    16'd48761,
    16'd48767,
    16'd48779,
    16'd48781,
    16'd48787,
    16'd48799,
    16'd48809,
    16'd48817,
    16'd48821,
    16'd48823,
    16'd48847,
    16'd48857,
    16'd48859,
    16'd48869,
    16'd48871,
    16'd48883,
    16'd48889,
    16'd48907,
    16'd48947,
    16'd48953,
    16'd48973,
    16'd48989,
    16'd48991,
    16'd49003,
    16'd49009,
    16'd49019,
    16'd49031,
    16'd49033,
    16'd49037,
    16'd49043,
    16'd49057,
    16'd49069,
    16'd49081,
    16'd49103,
    16'd49109,
    16'd49117,
    16'd49121,
    16'd49123,
    16'd49139,
    16'd49157,
    16'd49169,
    16'd49171,
    16'd49177,
    16'd49193,
    16'd49199,
    16'd49201,
    16'd49207,
    16'd49211,
    16'd49223,
    16'd49253,
    16'd49261,
    16'd49277,
    16'd49279,
    16'd49297,
    16'd49307,
    16'd49331,
    16'd49333,
    16'd49339,
    16'd49363,
    16'd49367,
    16'd49369,
    16'd49391,
    16'd49393,
    16'd49409,
    16'd49411,
    16'd49417,
    16'd49429,
    16'd49433,
    16'd49451,
    16'd49459,
    16'd49463,
    16'd49477,
    16'd49481,
    16'd49499,
    16'd49523,
    16'd49529,
    16'd49531,
    16'd49537,
    16'd49547,
    16'd49549,
    16'd49559,
    16'd49597,
    16'd49603,
    16'd49613,
    16'd49627,
    16'd49633,
    16'd49639,
    16'd49663,
    16'd49667,
    16'd49669,
    16'd49681,
    16'd49697,
    16'd49711,
    16'd49727,
    16'd49739,
    16'd49741,
    16'd49747,
    16'd49757,
    16'd49783,
    16'd49787,
    16'd49789,
    16'd49801,
    16'd49807,
    16'd49811,
    16'd49823,
    16'd49831,
    16'd49843,
    16'd49853,
    16'd49871,
    16'd49877,
    16'd49891,
    16'd49919,
    16'd49921,
    16'd49927,
    16'd49937,
    16'd49939,
    16'd49943,
    16'd49957,
    16'd49991,
    16'd49993,
    16'd49999,
    16'd50021,
    16'd50023,
    16'd50033,
    16'd50047,
    16'd50051,
    16'd50053,
    16'd50069,
    16'd50077,
    16'd50087,
    16'd50093,
    16'd50101,
    16'd50111,
    16'd50119,
    16'd50123,
    16'd50129,
    16'd50131,
    16'd50147,
    16'd50153,
    16'd50159,
    16'd50177,
    16'd50207,
    16'd50221,
    16'd50227,
    16'd50231,
    16'd50261,
    16'd50263,
    16'd50273,
    16'd50287,
    16'd50291,
    16'd50311,
    16'd50321,
    16'd50329,
    16'd50333,
    16'd50341,
    16'd50359,
    16'd50363,
    16'd50377,
    16'd50383,
    16'd50387,
    16'd50411,
    16'd50417,
    16'd50423,
    16'd50441,
    16'd50459,
    16'd50461,
    16'd50497,
    16'd50503,
    16'd50513,
    16'd50527,
    16'd50539,
    16'd50543,
    16'd50549,
    16'd50551,
    16'd50581,
    16'd50587,
    16'd50591,
    16'd50593,
    16'd50599,
    16'd50627,
    16'd50647,
    16'd50651,
    16'd50671,
    16'd50683,
    16'd50707,
    16'd50723,
    16'd50741,
    16'd50753,
    16'd50767,
    16'd50773,
    16'd50777,
    16'd50789,
    16'd50821,
    16'd50833,
    16'd50839,
    16'd50849,
    16'd50857,
    16'd50867,
    16'd50873,
    16'd50891,
    16'd50893,
    16'd50909,
    16'd50923,
    16'd50929,
    16'd50951,
    16'd50957,
    16'd50969,
    16'd50971,
    16'd50989,
    16'd50993,
    16'd51001,
    16'd51031,
    16'd51043,
    16'd51047,
    16'd51059,
    16'd51061,
    16'd51071,
    16'd51109,
    16'd51131,
    16'd51133,
    16'd51137,
    16'd51151,
    16'd51157,
    16'd51169,
    16'd51193,
    16'd51197,
    16'd51199,
    16'd51203,
    16'd51217,
    16'd51229,
    16'd51239,
    16'd51241,
    16'd51257,
    16'd51263,
    16'd51283,
    16'd51287,
    16'd51307,
    16'd51329,
    16'd51341,
    16'd51343,
    16'd51347,
    16'd51349,
    16'd51361,
    16'd51383,
    16'd51407,
    16'd51413,
    16'd51419,
    16'd51421,
    16'd51427,
    16'd51431,
    16'd51437,
    16'd51439,
    16'd51449,
    16'd51461,
    16'd51473,
    16'd51479,
    16'd51481,
    16'd51487,
    16'd51503,
    16'd51511,
    16'd51517,
    16'd51521,
    16'd51539,
    16'd51551,
    16'd51563,
    16'd51577,
    16'd51581,
    16'd51593,
    16'd51599,
    16'd51607,
    16'd51613,
    16'd51631,
    16'd51637,
    16'd51647,
    16'd51659,
    16'd51673,
    16'd51679,
    16'd51683,
    16'd51691,
    16'd51713,
    16'd51719,
    16'd51721,
    16'd51749,
    16'd51767,
    16'd51769,
    16'd51787,
    16'd51797,
    16'd51803,
    16'd51817,
    16'd51827,
    16'd51829,
    16'd51839,
    16'd51853,
    16'd51859,
    16'd51869,
    16'd51871,
    16'd51893,
    16'd51899,
    16'd51907,
    16'd51913,
    16'd51929,
    16'd51941,
    16'd51949,
    16'd51971,
    16'd51973,
    16'd51977,
    16'd51991,
    16'd52009,
    16'd52021,
    16'd52027,
    16'd52051,
    16'd52057,
    16'd52067,
    16'd52069,
    16'd52081,
    16'd52103,
    16'd52121,
    16'd52127,
    16'd52147,
    16'd52153,
    16'd52163,
    16'd52177,
    16'd52181,
    16'd52183,
    16'd52189,
    16'd52201,
    16'd52223,
    16'd52237,
    16'd52249,
    16'd52253,
    16'd52259,
    16'd52267,
    16'd52289,
    16'd52291,
    16'd52301,
    16'd52313,
    16'd52321,
    16'd52361,
    16'd52363,
    16'd52369,
    16'd52379,
    16'd52387,
    16'd52391,
    16'd52433,
    16'd52453,
    16'd52457,
    16'd52489,
    16'd52501,
    16'd52511,
    16'd52517,
    16'd52529,
    16'd52541,
    16'd52543,
    16'd52553,
    16'd52561,
    16'd52567,
    16'd52571,
    16'd52579,
    16'd52583,
    16'd52609,
    16'd52627,
    16'd52631,
    16'd52639,
    16'd52667,
    16'd52673,
    16'd52691,
    16'd52697,
    16'd52709,
    16'd52711,
    16'd52721,
    16'd52727,
    16'd52733,
    16'd52747,
    16'd52757,
    16'd52769,
    16'd52783,
    16'd52807,
    16'd52813,
    16'd52817,
    16'd52837,
    16'd52859,
    16'd52861,
    16'd52879,
    16'd52883,
    16'd52889,
    16'd52901,
    16'd52903,
    16'd52919,
    16'd52937,
    16'd52951,
    16'd52957,
    16'd52963,
    16'd52967,
    16'd52973,
    16'd52981,
    16'd52999,
    16'd53003,
    16'd53017,
    16'd53047,
    16'd53051,
    16'd53069,
    16'd53077,
    16'd53087,
    16'd53089,
    16'd53093,
    16'd53101,
    16'd53113,
    16'd53117,
    16'd53129,
    16'd53147,
    16'd53149,
    16'd53161,
    16'd53171,
    16'd53173,
    16'd53189,
    16'd53197,
    16'd53201,
    16'd53231,
    16'd53233,
    16'd53239,
    16'd53267,
    16'd53269,
    16'd53279,
    16'd53281,
    16'd53299,
    16'd53309,
    16'd53323,
    16'd53327,
    16'd53353,
    16'd53359,
    16'd53377,
    16'd53381,
    16'd53401,
    16'd53407,
    16'd53411,
    16'd53419,
    16'd53437,
    16'd53441,
    16'd53453,
    16'd53479,
    16'd53503,
    16'd53507,
    16'd53527,
    16'd53549,
    16'd53551,
    16'd53569,
    16'd53591,
    16'd53593,
    16'd53597,
    16'd53609,
    16'd53611,
    16'd53617,
    16'd53623,
    16'd53629,
    16'd53633,
    16'd53639,
    16'd53653,
    16'd53657,
    16'd53681,
    16'd53693,
    16'd53699,
    16'd53717,
    16'd53719,
    16'd53731,
    16'd53759,
    16'd53773,
    16'd53777,
    16'd53783,
    16'd53791,
    16'd53813,
    16'd53819,
    16'd53831,
    16'd53849,
    16'd53857,
    16'd53861,
    16'd53881,
    16'd53887,
    16'd53891,
    16'd53897,
    16'd53899,
    16'd53917,
    16'd53923,
    16'd53927,
    16'd53939,
    16'd53951,
    16'd53959,
    16'd53987,
    16'd53993,
    16'd54001,
    16'd54011,
    16'd54013,
    16'd54037,
    16'd54049,
    16'd54059,
    16'd54083,
    16'd54091,
    16'd54101,
    16'd54121,
    16'd54133,
    16'd54139,
    16'd54151,
    16'd54163,
    16'd54167,
    16'd54181,
    16'd54193,
    16'd54217,
    16'd54251,
    16'd54269,
    16'd54277,
    16'd54287,
    16'd54293,
    16'd54311,
    16'd54319,
    16'd54323,
    16'd54331,
    16'd54347,
    16'd54361,
    16'd54367,
    16'd54371,
    16'd54377,
    16'd54401,
    16'd54403,
    16'd54409,
    16'd54413,
    16'd54419,
    16'd54421,
    16'd54437,
    16'd54443,
    16'd54449,
    16'd54469,
    16'd54493,
    16'd54497,
    16'd54499,
    16'd54503,
    16'd54517,
    16'd54521,
    16'd54539,
    16'd54541,
    16'd54547,
    16'd54559,
    16'd54563,
    16'd54577,
    16'd54581,
    16'd54583,
    16'd54601,
    16'd54617,
    16'd54623,
    16'd54629,
    16'd54631,
    16'd54647,
    16'd54667,
    16'd54673,
    16'd54679,
    16'd54709,
    16'd54713,
    16'd54721,
    16'd54727,
    16'd54751,
    16'd54767,
    16'd54773,
    16'd54779,
    16'd54787,
    16'd54799,
    16'd54829,
    16'd54833,
    16'd54851,
    16'd54869,
    16'd54877,
    16'd54881,
    16'd54907,
    16'd54917,
    16'd54919,
    16'd54941,
    16'd54949,
    16'd54959,
    16'd54973,
    16'd54979,
    16'd54983,
    16'd55001,
    16'd55009,
    16'd55021,
    16'd55049,
    16'd55051,
    16'd55057,
    16'd55061,
    16'd55073,
    16'd55079,
    16'd55103,
    16'd55109,
    16'd55117,
    16'd55127,
    16'd55147,
    16'd55163,
    16'd55171,
    16'd55201,
    16'd55207,
    16'd55213,
    16'd55217,
    16'd55219,
    16'd55229,
    16'd55243,
    16'd55249,
    16'd55259,
    16'd55291,
    16'd55313,
    16'd55331,
    16'd55333,
    16'd55337,
    16'd55339,
    16'd55343,
    16'd55351,
    16'd55373,
    16'd55381,
    16'd55399,
    16'd55411,
    16'd55439,
    16'd55441,
    16'd55457,
    16'd55469,
    16'd55487,
    16'd55501,
    16'd55511,
    16'd55529,
    16'd55541,
    16'd55547,
    16'd55579,
    16'd55589,
    16'd55603,
    16'd55609,
    16'd55619,
    16'd55621,
    16'd55631,
    16'd55633,
    16'd55639,
    16'd55661,
    16'd55663,
    16'd55667,
    16'd55673,
    16'd55681,
    16'd55691,
    16'd55697,
    16'd55711,
    16'd55717,
    16'd55721,
    16'd55733,
    16'd55763,
    16'd55787,
    16'd55793,
    16'd55799,
    16'd55807,
    16'd55813,
    16'd55817,
    16'd55819,
    16'd55823,
    16'd55829,
    16'd55837,
    16'd55843,
    16'd55849,
    16'd55871,
    16'd55889,
    16'd55897,
    16'd55901,
    16'd55903,
    16'd55921,
    16'd55927,
    16'd55931,
    16'd55933,
    16'd55949,
    16'd55967,
    16'd55987,
    16'd55997,
    16'd56003,
    16'd56009,
    16'd56039,
    16'd56041,
    16'd56053,
    16'd56081,
    16'd56087,
    16'd56093,
    16'd56099,
    16'd56101,
    16'd56113,
    16'd56123,
    16'd56131,
    16'd56149,
    16'd56167,
    16'd56171,
    16'd56179,
    16'd56197,
    16'd56207,
    16'd56209,
    16'd56237,
    16'd56239,
    16'd56249,
    16'd56263,
    16'd56267,
    16'd56269,
    16'd56299,
    16'd56311,
    16'd56333,
    16'd56359,
    16'd56369,
    16'd56377,
    16'd56383,
    16'd56393,
    16'd56401,
    16'd56417,
    16'd56431,
    16'd56437,
    16'd56443,
    16'd56453,
    16'd56467,
    16'd56473,
    16'd56477,
    16'd56479,
    16'd56489,
    16'd56501,
    16'd56503,
    16'd56509,
    16'd56519,
    16'd56527,
    16'd56531,
    16'd56533,
    16'd56543,
    16'd56569,
    16'd56591,
    16'd56597,
    16'd56599,
    16'd56611,
    16'd56629,
    16'd56633,
    16'd56659,
    16'd56663,
    16'd56671,
    16'd56681,
    16'd56687,
    16'd56701,
    16'd56711,
    16'd56713,
    16'd56731,
    16'd56737,
    16'd56747,
    16'd56767,
    16'd56773,
    16'd56779,
    16'd56783,
    16'd56807,
    16'd56809,
    16'd56813,
    16'd56821,
    16'd56827,
    16'd56843,
    16'd56857,
    16'd56873,
    16'd56891,
    16'd56893,
    16'd56897,
    16'd56909,
    16'd56911,
    16'd56921,
    16'd56923,
    16'd56929,
    16'd56941,
    16'd56951,
    16'd56957,
    16'd56963,
    16'd56983,
    16'd56989,
    16'd56993,
    16'd56999,
    16'd57037,
    16'd57041,
    16'd57047,
    16'd57059,
    16'd57073,
    16'd57077,
    16'd57089,
    16'd57097,
    16'd57107,
    16'd57119,
    16'd57131,
    16'd57139,
    16'd57143,
    16'd57149,
    16'd57163,
    16'd57173,
    16'd57179,
    16'd57191,
    16'd57193,
    16'd57203,
    16'd57221,
    16'd57223,
    16'd57241,
    16'd57251,
    16'd57259,
    16'd57269,
    16'd57271,
    16'd57283,
    16'd57287,
    16'd57301,
    16'd57329,
    16'd57331,
    16'd57347,
    16'd57349,
    16'd57367,
    16'd57373,
    16'd57383,
    16'd57389,
    16'd57397,
    16'd57413,
    16'd57427,
    16'd57457,
    16'd57467,
    16'd57487,
    16'd57493,
    16'd57503,
    16'd57527,
    16'd57529,
    16'd57557,
    16'd57559,
    16'd57571,
    16'd57587,
    16'd57593,
    16'd57601,
    16'd57637,
    16'd57641,
    16'd57649,
    16'd57653,
    16'd57667,
    16'd57679,
    16'd57689,
    16'd57697,
    16'd57709,
    16'd57713,
    16'd57719,
    16'd57727,
    16'd57731,
    16'd57737,
    16'd57751,
    16'd57773,
    16'd57781,
    16'd57787,
    16'd57791,
    16'd57793,
    16'd57803,
    16'd57809,
    16'd57829,
    16'd57839,
    16'd57847,
    16'd57853,
    16'd57859,
    16'd57881,
    16'd57899,
    16'd57901,
    16'd57917,
    16'd57923,
    16'd57943,
    16'd57947,
    16'd57973,
    16'd57977,
    16'd57991,
    16'd58013,
    16'd58027,
    16'd58031,
    16'd58043,
    16'd58049,
    16'd58057,
    16'd58061,
    16'd58067,
    16'd58073,
    16'd58099,
    16'd58109,
    16'd58111,
    16'd58129,
    16'd58147,
    16'd58151,
    16'd58153,
    16'd58169,
    16'd58171,
    16'd58189,
    16'd58193,
    16'd58199,
    16'd58207,
    16'd58211,
    16'd58217,
    16'd58229,
    16'd58231,
    16'd58237,
    16'd58243,
    16'd58271,
    16'd58309,
    16'd58313,
    16'd58321,
    16'd58337,
    16'd58363,
    16'd58367,
    16'd58369,
    16'd58379,
    16'd58391,
    16'd58393,
    16'd58403,
    16'd58411,
    16'd58417,
    16'd58427,
    16'd58439,
    16'd58441,
    16'd58451,
    16'd58453,
    16'd58477,
    16'd58481,
    16'd58511,
    16'd58537,
    16'd58543,
    16'd58549,
    16'd58567,
    16'd58573,
    16'd58579,
    16'd58601,
    16'd58603,
    16'd58613,
    16'd58631,
    16'd58657,
    16'd58661,
    16'd58679,
    16'd58687,
    16'd58693,
    16'd58699,
    16'd58711,
    16'd58727,
    16'd58733,
    16'd58741,
    16'd58757,
    16'd58763,
    16'd58771,
    16'd58787,
    16'd58789,
    16'd58831,
    16'd58889,
    16'd58897,
    16'd58901,
    16'd58907,
    16'd58909,
    16'd58913,
    16'd58921,
    16'd58937,
    16'd58943,
    16'd58963,
    16'd58967,
    16'd58979,
    16'd58991,
    16'd58997,
    16'd59009,
    16'd59011,
    16'd59021,
    16'd59023,
    16'd59029,
    16'd59051,
    16'd59053,
    16'd59063,
    16'd59069,
    16'd59077,
    16'd59083,
    16'd59093,
    16'd59107,
    16'd59113,
    16'd59119,
    16'd59123,
    16'd59141,
    16'd59149,
    16'd59159,
    16'd59167,
    16'd59183,
    16'd59197,
    16'd59207,
    16'd59209,
    16'd59219,
    16'd59221,
    16'd59233,
    16'd59239,
    16'd59243,
    16'd59263,
    16'd59273,
    16'd59281,
    16'd59333,
    16'd59341,
    16'd59351,
    16'd59357,
    16'd59359,
    16'd59369,
    16'd59377,
    16'd59387,
    16'd59393,
    16'd59399,
    16'd59407,
    16'd59417,
    16'd59419,
    16'd59441,
    16'd59443,
    16'd59447,
    16'd59453,
    16'd59467,
    16'd59471,
    16'd59473,
    16'd59497,
    16'd59509,
    16'd59513,
    16'd59539,
    16'd59557,
    16'd59561,
    16'd59567,
    16'd59581,
    16'd59611,
    16'd59617,
    16'd59621,
    16'd59627,
    16'd59629,
    16'd59651,
    16'd59659,
    16'd59663,
    16'd59669,
    16'd59671,
    16'd59693,
    16'd59699,
    16'd59707,
    16'd59723,
    16'd59729,
    16'd59743,
    16'd59747,
    16'd59753,
    16'd59771,
    16'd59779,
    16'd59791,
    16'd59797,
    16'd59809,
    16'd59833,
    16'd59863,
    16'd59879,
    16'd59887,
    16'd59921,
    16'd59929,
    16'd59951,
    16'd59957,
    16'd59971,
    16'd59981,
    16'd59999,
    16'd60013,
    16'd60017,
    16'd60029,
    16'd60037,
    16'd60041,
    16'd60077,
    16'd60083,
    16'd60089,
    16'd60091,
    16'd60101,
    16'd60103,
    16'd60107,
    16'd60127,
    16'd60133,
    16'd60139,
    16'd60149,
    16'd60161,
    16'd60167,
    16'd60169,
    16'd60209,
    16'd60217,
    16'd60223,
    16'd60251,
    16'd60257,
    16'd60259,
    16'd60271,
    16'd60289,
    16'd60293,
    16'd60317,
    16'd60331,
    16'd60337,
    16'd60343,
    16'd60353,
    16'd60373,
    16'd60383,
    16'd60397,
    16'd60413,
    16'd60427,
    16'd60443,
    16'd60449,
    16'd60457,
    16'd60493,
    16'd60497,
    16'd60509,
    16'd60521,
    16'd60527,
    16'd60539,
    16'd60589,
    16'd60601,
    16'd60607,
    16'd60611,
    16'd60617,
    16'd60623,
    16'd60631,
    16'd60637,
    16'd60647,
    16'd60649,
    16'd60659,
    16'd60661,
    16'd60679,
    16'd60689,
    16'd60703,
    16'd60719,
    16'd60727,
    16'd60733,
    16'd60737,
    16'd60757,
    16'd60761,
    16'd60763,
    16'd60773,
    16'd60779,
    16'd60793,
    16'd60811,
    16'd60821,
    16'd60859,
    16'd60869,
    16'd60887,
    16'd60889,
    16'd60899,
    16'd60901,
    16'd60913,
    16'd60917,
    16'd60919,
    16'd60923,
    16'd60937,
    16'd60943,
    16'd60953,
    16'd60961,
    16'd61001,
    16'd61007,
    16'd61027,
    16'd61031,
    16'd61043,
    16'd61051,
    16'd61057,
    16'd61091,
    16'd61099,
    16'd61121,
    16'd61129,
    16'd61141,
    16'd61151,
    16'd61153,
    16'd61169,
    16'd61211,
    16'd61223,
    16'd61231,
    16'd61253,
    16'd61261,
    16'd61283,
    16'd61291,
    16'd61297,
    16'd61331,
    16'd61333,
    16'd61339,
    16'd61343,
    16'd61357,
    16'd61363,
    16'd61379,
    16'd61381,
    16'd61403,
    16'd61409,
    16'd61417,
    16'd61441,
    16'd61463,
    16'd61469,
    16'd61471,
    16'd61483,
    16'd61487,
    16'd61493,
    16'd61507,
    16'd61511,
    16'd61519,
    16'd61543,
    16'd61547,
    16'd61553,
    16'd61559,
    16'd61561,
    16'd61583,
    16'd61603,
    16'd61609,
    16'd61613,
    16'd61627,
    16'd61631,
    16'd61637,
    16'd61643,
    16'd61651,
    16'd61657,
    16'd61667,
    16'd61673,
    16'd61681,
    16'd61687,
    16'd61703,
    16'd61717,
    16'd61723,
    16'd61729,
    16'd61751,
    16'd61757,
    16'd61781,
    16'd61813,
    16'd61819,
    16'd61837,
    16'd61843,
    16'd61861,
    16'd61871,
    16'd61879,
    16'd61909,
    16'd61927,
    16'd61933,
    16'd61949,
    16'd61961,
    16'd61967,
    16'd61979,
    16'd61981,
    16'd61987,
    16'd61991,
    16'd62003,
    16'd62011,
    16'd62017,
    16'd62039,
    16'd62047,
    16'd62053,
    16'd62057,
    16'd62071,
    16'd62081,
    16'd62099,
    16'd62119,
    16'd62129,
    16'd62131,
    16'd62137,
    16'd62141,
    16'd62143,
    16'd62171,
    16'd62189,
    16'd62191,
    16'd62201,
    16'd62207,
    16'd62213,
    16'd62219,
    16'd62233,
    16'd62273,
    16'd62297,
    16'd62299,
    16'd62303,
    16'd62311,
    16'd62323,
    16'd62327,
    16'd62347,
    16'd62351,
    16'd62383,
    16'd62401,
    16'd62417,
    16'd62423,
    16'd62459,
    16'd62467,
    16'd62473,
    16'd62477,
    16'd62483,
    16'd62497,
    16'd62501,
    16'd62507,
    16'd62533,
    16'd62539,
    16'd62549,
    16'd62563,
    16'd62581,
    16'd62591,
    16'd62597,
    16'd62603,
    16'd62617,
    16'd62627,
    16'd62633,
    16'd62639,
    16'd62653,
    16'd62659,
    16'd62683,
    16'd62687,
    16'd62701,
    16'd62723,
    16'd62731,
    16'd62743,
    16'd62753,
    16'd62761,
    16'd62773,
    16'd62791,
    16'd62801,
    16'd62819,
    16'd62827,
    16'd62851,
    16'd62861,
    16'd62869,
    16'd62873,
    16'd62897,
    16'd62903,
    16'd62921,
    16'd62927,
    16'd62929,
    16'd62939,
    16'd62969,
    16'd62971,
    16'd62981,
    16'd62983,
    16'd62987,
    16'd62989,
    16'd63029,
    16'd63031,
    16'd63059,
    16'd63067,
    16'd63073,
    16'd63079,
    16'd63097,
    16'd63103,
    16'd63113,
    16'd63127,
    16'd63131,
    16'd63149,
    16'd63179,
    16'd63197,
    16'd63199,
    16'd63211,
    16'd63241,
    16'd63247,
    16'd63277,
    16'd63281,
    16'd63299,
    16'd63311,
    16'd63313,
    16'd63317,
    16'd63331,
    16'd63337,
    16'd63347,
    16'd63353,
    16'd63361,
    16'd63367,
    16'd63377,
    16'd63389,
    16'd63391,
    16'd63397,
    16'd63409,
    16'd63419,
    16'd63421,
    16'd63439,
    16'd63443,
    16'd63463,
    16'd63467,
    16'd63473,
    16'd63487,
    16'd63493,
    16'd63499,
    16'd63521,
    16'd63527,
    16'd63533,
    16'd63541,
    16'd63559,
    16'd63577,
    16'd63587,
    16'd63589,
    16'd63599,
    16'd63601,
    16'd63607,
    16'd63611,
    16'd63617,
    16'd63629,
    16'd63647,
    16'd63649,
    16'd63659,
    16'd63667,
    16'd63671,
    16'd63689,
    16'd63691,
    16'd63697,
    16'd63703,
    16'd63709,
    16'd63719,
    16'd63727,
    16'd63737,
    16'd63743,
    16'd63761,
    16'd63773,
    16'd63781,
    16'd63793,
    16'd63799,
    16'd63803,
    16'd63809,
    16'd63823,
    16'd63839,
    16'd63841,
    16'd63853,
    16'd63857,
    16'd63863,
    16'd63901,
    16'd63907,
    16'd63913,
    16'd63929,
    16'd63949,
    16'd63977,
    16'd63997,
    16'd64007,
    16'd64013,
    16'd64019,
    16'd64033,
    16'd64037,
    16'd64063,
    16'd64067,
    16'd64081,
    16'd64091,
    16'd64109,
    16'd64123,
    16'd64151,
    16'd64153,
    16'd64157,
    16'd64171,
    16'd64187,
    16'd64189,
    16'd64217,
    16'd64223,
    16'd64231,
    16'd64237,
    16'd64271,
    16'd64279,
    16'd64283,
    16'd64301,
    16'd64303,
    16'd64319,
    16'd64327,
    16'd64333,
    16'd64373,
    16'd64381,
    16'd64399,
    16'd64403,
    16'd64433,
    16'd64439,
    16'd64451,
    16'd64453,
    16'd64483,
    16'd64489,
    16'd64499,
    16'd64513,
    16'd64553,
    16'd64567,
    16'd64577,
    16'd64579,
    16'd64591,
    16'd64601,
    16'd64609,
    16'd64613,
    16'd64621,
    16'd64627,
    16'd64633,
    16'd64661,
    16'd64663,
    16'd64667,
    16'd64679,
    16'd64693,
    16'd64709,
    16'd64717,
    16'd64747,
    16'd64763,
    16'd64781,
    16'd64783,
    16'd64793,
    16'd64811,
    16'd64817,
    16'd64849,
    16'd64853,
    16'd64871,
    16'd64877,
    16'd64879,
    16'd64891,
    16'd64901,
    16'd64919,
    16'd64921,
    16'd64927,
    16'd64937,
    16'd64951,
    16'd64969,
    16'd64997,
    16'd65003,
    16'd65011,
    16'd65027,
    16'd65029,
    16'd65033,
    16'd65053,
    16'd65063,
    16'd65071,
    16'd65089,
    16'd65099,
    16'd65101,
    16'd65111,
    16'd65119,
    16'd65123,
    16'd65129,
    16'd65141,
    16'd65147,
    16'd65167,
    16'd65171,
    16'd65173,
    16'd65179,
    16'd65183,
    16'd65203,
    16'd65213,
    16'd65239,
    16'd65257,
    16'd65267,
    16'd65269,
    16'd65287,
    16'd65293,
    16'd65309,
    16'd65323,
    16'd65327,
    16'd65353,
    16'd65357,
    16'd65371,
    16'd65381,
    16'd65393,
    16'd65407,
    16'd65413,
    16'd65419,
    16'd65423,
    16'd65437,
    16'd65447,
    16'd65449,
    16'd65479,
    16'd65497,
    16'd65519,
    16'd65521
};

parameter IDLE = 0;
parameter CALC = 1;

// wire [15:0] test;
// assign test = PrimeArray[16*3 +: 16];

// ========== reg and wire =========
reg  [       15:0] low, low_nxt;
reg  [       15:0] mid, mid_nxt;
reg  [       15:0] high, high_nxt;
reg  [  WIDTH-1:0] num_reg;
reg  [        2:0] state, state_nxt;

reg                finish_nxt;
reg                IsPrime_nxt;

wire [       15:0] CurrentEntry;
// wire [       15:0] cool;

assign CurrentEntry = PrimeArray[16*(mid-1) +: 16];
// assign cool = PrimeArray[0: 15];

// reg AssumePrime;

// ========== Combinational =========
// state
always @(*) begin
    state_nxt = state;
    if (state == IDLE) begin
        if (start) state_nxt = CALC;
    end else begin
        // hit
        if (num_reg == CurrentEntry) begin
            state_nxt = IDLE;
        end else if (low >= high) begin // search not found
            state_nxt = IDLE;
        end
    end
end

// finish and IsPrime
always @(*) begin
    finish_nxt = 0;
    IsPrime_nxt = 0;
    if (state == CALC) begin
        // hit
        if (num_reg == CurrentEntry) begin
            finish_nxt = 1;
            IsPrime_nxt = 1;
        end else if (low >= high) begin // search not found
            finish_nxt = 1;
            IsPrime_nxt = 0;
        end
    end
end

// low_nxt, mid_nxt, high_nxt
always @(*) begin
    low_nxt  = low;
    mid_nxt  = mid;
    high_nxt = high;
    if (state == CALC) begin
        if (num_reg < CurrentEntry) begin
            high_nxt = mid - 1;
            mid_nxt  = (low + (mid-1)) >> 1;
        end else if (num_reg > CurrentEntry) begin
            low_nxt = mid + 1;
            mid_nxt = ((mid+1) + high) >> 1;
        end
    end
end

// ========== Sequential =========
// state
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
    end else begin
        state <= state_nxt;
    end
end

// num_reg
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        num_reg <= 0;
    end else begin
        if (start) begin
            num_reg <= num;
        end else begin
            num_reg <= num_reg;
        end
    end
end

// binary search index
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        low  <= 1;
        mid  <= (PRIME_COUNT) >> 1;
        high <= (PRIME_COUNT);
    end else begin
        low  <= low_nxt;
        mid  <= mid_nxt;
        high <= high_nxt;
    end
end

// output
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        finish  <= 0;
        IsPrime <= 0;
    end else begin
        finish  <= finish_nxt;
        IsPrime <= IsPrime_nxt;
    end
end

// AssumePrime
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        AssumePrime <= 1;
    end else begin
        if (finish && !IsPrime) begin
            AssumePrime <= 0;
        end
        else begin
            AssumePrime <= AssumePrime;
        end
    end
end

endmodule