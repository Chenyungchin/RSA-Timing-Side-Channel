module add(
    input [255:0] a,
    input [255:0] b,
    output [255:0] c
);
    assign c = a + b;

endmodule