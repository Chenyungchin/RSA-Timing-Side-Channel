module CheckPrime_comb #(parameter WIDTH = 8) (
    // input
    input      [  WIDTH-1:0] num,
    // output
    output reg               AssumePrime
);
// assign test = PrimeArray[16*3 +: 16];

always @(*) begin
    AssumePrime = 0;
	if (num==16'd2) begin
		AssumePrime = 1;
	end	else if (num==16'd3) begin
		AssumePrime = 1;
	end	else if (num==16'd5) begin
		AssumePrime = 1;
	end	else if (num==16'd7) begin
		AssumePrime = 1;
	end	else if (num==16'd11) begin
		AssumePrime = 1;
	end	else if (num==16'd13) begin
		AssumePrime = 1;
	end	else if (num==16'd17) begin
		AssumePrime = 1;
	end	else if (num==16'd19) begin
		AssumePrime = 1;
	end	else if (num==16'd23) begin
		AssumePrime = 1;
	end	else if (num==16'd29) begin
		AssumePrime = 1;
	end	else if (num==16'd31) begin
		AssumePrime = 1;
	end	else if (num==16'd37) begin
		AssumePrime = 1;
	end	else if (num==16'd41) begin
		AssumePrime = 1;
	end	else if (num==16'd43) begin
		AssumePrime = 1;
	end	else if (num==16'd47) begin
		AssumePrime = 1;
	end	else if (num==16'd53) begin
		AssumePrime = 1;
	end	else if (num==16'd59) begin
		AssumePrime = 1;
	end	else if (num==16'd61) begin
		AssumePrime = 1;
	end	else if (num==16'd67) begin
		AssumePrime = 1;
	end	else if (num==16'd71) begin
		AssumePrime = 1;
	end	else if (num==16'd73) begin
		AssumePrime = 1;
	end	else if (num==16'd79) begin
		AssumePrime = 1;
	end	else if (num==16'd83) begin
		AssumePrime = 1;
	end	else if (num==16'd89) begin
		AssumePrime = 1;
	end	else if (num==16'd97) begin
		AssumePrime = 1;
	end	else if (num==16'd101) begin
		AssumePrime = 1;
	end	else if (num==16'd103) begin
		AssumePrime = 1;
	end	else if (num==16'd107) begin
		AssumePrime = 1;
	end	else if (num==16'd109) begin
		AssumePrime = 1;
	end	else if (num==16'd113) begin
		AssumePrime = 1;
	end	else if (num==16'd127) begin
		AssumePrime = 1;
	end	else if (num==16'd131) begin
		AssumePrime = 1;
	end	else if (num==16'd137) begin
		AssumePrime = 1;
	end	else if (num==16'd139) begin
		AssumePrime = 1;
	end	else if (num==16'd149) begin
		AssumePrime = 1;
	end	else if (num==16'd151) begin
		AssumePrime = 1;
	end	else if (num==16'd157) begin
		AssumePrime = 1;
	end	else if (num==16'd163) begin
		AssumePrime = 1;
	end	else if (num==16'd167) begin
		AssumePrime = 1;
	end	else if (num==16'd173) begin
		AssumePrime = 1;
	end	else if (num==16'd179) begin
		AssumePrime = 1;
	end	else if (num==16'd181) begin
		AssumePrime = 1;
	end	else if (num==16'd191) begin
		AssumePrime = 1;
	end	else if (num==16'd193) begin
		AssumePrime = 1;
	end	else if (num==16'd197) begin
		AssumePrime = 1;
	end	else if (num==16'd199) begin
		AssumePrime = 1;
	end	else if (num==16'd211) begin
		AssumePrime = 1;
	end	else if (num==16'd223) begin
		AssumePrime = 1;
	end	else if (num==16'd227) begin
		AssumePrime = 1;
	end	else if (num==16'd229) begin
		AssumePrime = 1;
	end	else if (num==16'd233) begin
		AssumePrime = 1;
	end	else if (num==16'd239) begin
		AssumePrime = 1;
	end	else if (num==16'd241) begin
		AssumePrime = 1;
	end	else if (num==16'd251) begin
		AssumePrime = 1;
	end	else if (num==16'd257) begin
		AssumePrime = 1;
	end	else if (num==16'd263) begin
		AssumePrime = 1;
	end	else if (num==16'd269) begin
		AssumePrime = 1;
	end	else if (num==16'd271) begin
		AssumePrime = 1;
	end	else if (num==16'd277) begin
		AssumePrime = 1;
	end	else if (num==16'd281) begin
		AssumePrime = 1;
	end	else if (num==16'd283) begin
		AssumePrime = 1;
	end	else if (num==16'd293) begin
		AssumePrime = 1;
	end	else if (num==16'd307) begin
		AssumePrime = 1;
	end	else if (num==16'd311) begin
		AssumePrime = 1;
	end	else if (num==16'd313) begin
		AssumePrime = 1;
	end	else if (num==16'd317) begin
		AssumePrime = 1;
	end	else if (num==16'd331) begin
		AssumePrime = 1;
	end	else if (num==16'd337) begin
		AssumePrime = 1;
	end	else if (num==16'd347) begin
		AssumePrime = 1;
	end	else if (num==16'd349) begin
		AssumePrime = 1;
	end	else if (num==16'd353) begin
		AssumePrime = 1;
	end	else if (num==16'd359) begin
		AssumePrime = 1;
	end	else if (num==16'd367) begin
		AssumePrime = 1;
	end	else if (num==16'd373) begin
		AssumePrime = 1;
	end	else if (num==16'd379) begin
		AssumePrime = 1;
	end	else if (num==16'd383) begin
		AssumePrime = 1;
	end	else if (num==16'd389) begin
		AssumePrime = 1;
	end	else if (num==16'd397) begin
		AssumePrime = 1;
	end	else if (num==16'd401) begin
		AssumePrime = 1;
	end	else if (num==16'd409) begin
		AssumePrime = 1;
	end	else if (num==16'd419) begin
		AssumePrime = 1;
	end	else if (num==16'd421) begin
		AssumePrime = 1;
	end	else if (num==16'd431) begin
		AssumePrime = 1;
	end	else if (num==16'd433) begin
		AssumePrime = 1;
	end	else if (num==16'd439) begin
		AssumePrime = 1;
	end	else if (num==16'd443) begin
		AssumePrime = 1;
	end	else if (num==16'd449) begin
		AssumePrime = 1;
	end	else if (num==16'd457) begin
		AssumePrime = 1;
	end	else if (num==16'd461) begin
		AssumePrime = 1;
	end	else if (num==16'd463) begin
		AssumePrime = 1;
	end	else if (num==16'd467) begin
		AssumePrime = 1;
	end	else if (num==16'd479) begin
		AssumePrime = 1;
	end	else if (num==16'd487) begin
		AssumePrime = 1;
	end	else if (num==16'd491) begin
		AssumePrime = 1;
	end	else if (num==16'd499) begin
		AssumePrime = 1;
	end	else if (num==16'd503) begin
		AssumePrime = 1;
	end	else if (num==16'd509) begin
		AssumePrime = 1;
	end	else if (num==16'd521) begin
		AssumePrime = 1;
	end	else if (num==16'd523) begin
		AssumePrime = 1;
	end	else if (num==16'd541) begin
		AssumePrime = 1;
	end	else if (num==16'd547) begin
		AssumePrime = 1;
	end	else if (num==16'd557) begin
		AssumePrime = 1;
	end	else if (num==16'd563) begin
		AssumePrime = 1;
	end	else if (num==16'd569) begin
		AssumePrime = 1;
	end	else if (num==16'd571) begin
		AssumePrime = 1;
	end	else if (num==16'd577) begin
		AssumePrime = 1;
	end	else if (num==16'd587) begin
		AssumePrime = 1;
	end	else if (num==16'd593) begin
		AssumePrime = 1;
	end	else if (num==16'd599) begin
		AssumePrime = 1;
	end	else if (num==16'd601) begin
		AssumePrime = 1;
	end	else if (num==16'd607) begin
		AssumePrime = 1;
	end	else if (num==16'd613) begin
		AssumePrime = 1;
	end	else if (num==16'd617) begin
		AssumePrime = 1;
	end	else if (num==16'd619) begin
		AssumePrime = 1;
	end	else if (num==16'd631) begin
		AssumePrime = 1;
	end	else if (num==16'd641) begin
		AssumePrime = 1;
	end	else if (num==16'd643) begin
		AssumePrime = 1;
	end	else if (num==16'd647) begin
		AssumePrime = 1;
	end	else if (num==16'd653) begin
		AssumePrime = 1;
	end	else if (num==16'd659) begin
		AssumePrime = 1;
	end	else if (num==16'd661) begin
		AssumePrime = 1;
	end	else if (num==16'd673) begin
		AssumePrime = 1;
	end	else if (num==16'd677) begin
		AssumePrime = 1;
	end	else if (num==16'd683) begin
		AssumePrime = 1;
	end	else if (num==16'd691) begin
		AssumePrime = 1;
	end	else if (num==16'd701) begin
		AssumePrime = 1;
	end	else if (num==16'd709) begin
		AssumePrime = 1;
	end	else if (num==16'd719) begin
		AssumePrime = 1;
	end	else if (num==16'd727) begin
		AssumePrime = 1;
	end	else if (num==16'd733) begin
		AssumePrime = 1;
	end	else if (num==16'd739) begin
		AssumePrime = 1;
	end	else if (num==16'd743) begin
		AssumePrime = 1;
	end	else if (num==16'd751) begin
		AssumePrime = 1;
	end	else if (num==16'd757) begin
		AssumePrime = 1;
	end	else if (num==16'd761) begin
		AssumePrime = 1;
	end	else if (num==16'd769) begin
		AssumePrime = 1;
	end	else if (num==16'd773) begin
		AssumePrime = 1;
	end	else if (num==16'd787) begin
		AssumePrime = 1;
	end	else if (num==16'd797) begin
		AssumePrime = 1;
	end	else if (num==16'd809) begin
		AssumePrime = 1;
	end	else if (num==16'd811) begin
		AssumePrime = 1;
	end	else if (num==16'd821) begin
		AssumePrime = 1;
	end	else if (num==16'd823) begin
		AssumePrime = 1;
	end	else if (num==16'd827) begin
		AssumePrime = 1;
	end	else if (num==16'd829) begin
		AssumePrime = 1;
	end	else if (num==16'd839) begin
		AssumePrime = 1;
	end	else if (num==16'd853) begin
		AssumePrime = 1;
	end	else if (num==16'd857) begin
		AssumePrime = 1;
	end	else if (num==16'd859) begin
		AssumePrime = 1;
	end	else if (num==16'd863) begin
		AssumePrime = 1;
	end	else if (num==16'd877) begin
		AssumePrime = 1;
	end	else if (num==16'd881) begin
		AssumePrime = 1;
	end	else if (num==16'd883) begin
		AssumePrime = 1;
	end	else if (num==16'd887) begin
		AssumePrime = 1;
	end	else if (num==16'd907) begin
		AssumePrime = 1;
	end	else if (num==16'd911) begin
		AssumePrime = 1;
	end	else if (num==16'd919) begin
		AssumePrime = 1;
	end	else if (num==16'd929) begin
		AssumePrime = 1;
	end	else if (num==16'd937) begin
		AssumePrime = 1;
	end	else if (num==16'd941) begin
		AssumePrime = 1;
	end	else if (num==16'd947) begin
		AssumePrime = 1;
	end	else if (num==16'd953) begin
		AssumePrime = 1;
	end	else if (num==16'd967) begin
		AssumePrime = 1;
	end	else if (num==16'd971) begin
		AssumePrime = 1;
	end	else if (num==16'd977) begin
		AssumePrime = 1;
	end	else if (num==16'd983) begin
		AssumePrime = 1;
	end	else if (num==16'd991) begin
		AssumePrime = 1;
	end	else if (num==16'd997) begin
		AssumePrime = 1;
	end	else if (num==16'd1009) begin
		AssumePrime = 1;
	end	else if (num==16'd1013) begin
		AssumePrime = 1;
	end	else if (num==16'd1019) begin
		AssumePrime = 1;
	end	else if (num==16'd1021) begin
		AssumePrime = 1;
	end	else if (num==16'd1031) begin
		AssumePrime = 1;
	end	else if (num==16'd1033) begin
		AssumePrime = 1;
	end	else if (num==16'd1039) begin
		AssumePrime = 1;
	end	else if (num==16'd1049) begin
		AssumePrime = 1;
	end	else if (num==16'd1051) begin
		AssumePrime = 1;
	end	else if (num==16'd1061) begin
		AssumePrime = 1;
	end	else if (num==16'd1063) begin
		AssumePrime = 1;
	end	else if (num==16'd1069) begin
		AssumePrime = 1;
	end	else if (num==16'd1087) begin
		AssumePrime = 1;
	end	else if (num==16'd1091) begin
		AssumePrime = 1;
	end	else if (num==16'd1093) begin
		AssumePrime = 1;
	end	else if (num==16'd1097) begin
		AssumePrime = 1;
	end	else if (num==16'd1103) begin
		AssumePrime = 1;
	end	else if (num==16'd1109) begin
		AssumePrime = 1;
	end	else if (num==16'd1117) begin
		AssumePrime = 1;
	end	else if (num==16'd1123) begin
		AssumePrime = 1;
	end	else if (num==16'd1129) begin
		AssumePrime = 1;
	end	else if (num==16'd1151) begin
		AssumePrime = 1;
	end	else if (num==16'd1153) begin
		AssumePrime = 1;
	end	else if (num==16'd1163) begin
		AssumePrime = 1;
	end	else if (num==16'd1171) begin
		AssumePrime = 1;
	end	else if (num==16'd1181) begin
		AssumePrime = 1;
	end	else if (num==16'd1187) begin
		AssumePrime = 1;
	end	else if (num==16'd1193) begin
		AssumePrime = 1;
	end	else if (num==16'd1201) begin
		AssumePrime = 1;
	end	else if (num==16'd1213) begin
		AssumePrime = 1;
	end	else if (num==16'd1217) begin
		AssumePrime = 1;
	end	else if (num==16'd1223) begin
		AssumePrime = 1;
	end	else if (num==16'd1229) begin
		AssumePrime = 1;
	end	else if (num==16'd1231) begin
		AssumePrime = 1;
	end	else if (num==16'd1237) begin
		AssumePrime = 1;
	end	else if (num==16'd1249) begin
		AssumePrime = 1;
	end	else if (num==16'd1259) begin
		AssumePrime = 1;
	end	else if (num==16'd1277) begin
		AssumePrime = 1;
	end	else if (num==16'd1279) begin
		AssumePrime = 1;
	end	else if (num==16'd1283) begin
		AssumePrime = 1;
	end	else if (num==16'd1289) begin
		AssumePrime = 1;
	end	else if (num==16'd1291) begin
		AssumePrime = 1;
	end	else if (num==16'd1297) begin
		AssumePrime = 1;
	end	else if (num==16'd1301) begin
		AssumePrime = 1;
	end	else if (num==16'd1303) begin
		AssumePrime = 1;
	end	else if (num==16'd1307) begin
		AssumePrime = 1;
	end	else if (num==16'd1319) begin
		AssumePrime = 1;
	end	else if (num==16'd1321) begin
		AssumePrime = 1;
	end	else if (num==16'd1327) begin
		AssumePrime = 1;
	end	else if (num==16'd1361) begin
		AssumePrime = 1;
	end	else if (num==16'd1367) begin
		AssumePrime = 1;
	end	else if (num==16'd1373) begin
		AssumePrime = 1;
	end	else if (num==16'd1381) begin
		AssumePrime = 1;
	end	else if (num==16'd1399) begin
		AssumePrime = 1;
	end	else if (num==16'd1409) begin
		AssumePrime = 1;
	end	else if (num==16'd1423) begin
		AssumePrime = 1;
	end	else if (num==16'd1427) begin
		AssumePrime = 1;
	end	else if (num==16'd1429) begin
		AssumePrime = 1;
	end	else if (num==16'd1433) begin
		AssumePrime = 1;
	end	else if (num==16'd1439) begin
		AssumePrime = 1;
	end	else if (num==16'd1447) begin
		AssumePrime = 1;
	end	else if (num==16'd1451) begin
		AssumePrime = 1;
	end	else if (num==16'd1453) begin
		AssumePrime = 1;
	end	else if (num==16'd1459) begin
		AssumePrime = 1;
	end	else if (num==16'd1471) begin
		AssumePrime = 1;
	end	else if (num==16'd1481) begin
		AssumePrime = 1;
	end	else if (num==16'd1483) begin
		AssumePrime = 1;
	end	else if (num==16'd1487) begin
		AssumePrime = 1;
	end	else if (num==16'd1489) begin
		AssumePrime = 1;
	end	else if (num==16'd1493) begin
		AssumePrime = 1;
	end	else if (num==16'd1499) begin
		AssumePrime = 1;
	end	else if (num==16'd1511) begin
		AssumePrime = 1;
	end	else if (num==16'd1523) begin
		AssumePrime = 1;
	end	else if (num==16'd1531) begin
		AssumePrime = 1;
	end	else if (num==16'd1543) begin
		AssumePrime = 1;
	end	else if (num==16'd1549) begin
		AssumePrime = 1;
	end	else if (num==16'd1553) begin
		AssumePrime = 1;
	end	else if (num==16'd1559) begin
		AssumePrime = 1;
	end	else if (num==16'd1567) begin
		AssumePrime = 1;
	end	else if (num==16'd1571) begin
		AssumePrime = 1;
	end	else if (num==16'd1579) begin
		AssumePrime = 1;
	end	else if (num==16'd1583) begin
		AssumePrime = 1;
	end	else if (num==16'd1597) begin
		AssumePrime = 1;
	end	else if (num==16'd1601) begin
		AssumePrime = 1;
	end	else if (num==16'd1607) begin
		AssumePrime = 1;
	end	else if (num==16'd1609) begin
		AssumePrime = 1;
	end	else if (num==16'd1613) begin
		AssumePrime = 1;
	end	else if (num==16'd1619) begin
		AssumePrime = 1;
	end	else if (num==16'd1621) begin
		AssumePrime = 1;
	end	else if (num==16'd1627) begin
		AssumePrime = 1;
	end	else if (num==16'd1637) begin
		AssumePrime = 1;
	end	else if (num==16'd1657) begin
		AssumePrime = 1;
	end	else if (num==16'd1663) begin
		AssumePrime = 1;
	end	else if (num==16'd1667) begin
		AssumePrime = 1;
	end	else if (num==16'd1669) begin
		AssumePrime = 1;
	end	else if (num==16'd1693) begin
		AssumePrime = 1;
	end	else if (num==16'd1697) begin
		AssumePrime = 1;
	end	else if (num==16'd1699) begin
		AssumePrime = 1;
	end	else if (num==16'd1709) begin
		AssumePrime = 1;
	end	else if (num==16'd1721) begin
		AssumePrime = 1;
	end	else if (num==16'd1723) begin
		AssumePrime = 1;
	end	else if (num==16'd1733) begin
		AssumePrime = 1;
	end	else if (num==16'd1741) begin
		AssumePrime = 1;
	end	else if (num==16'd1747) begin
		AssumePrime = 1;
	end	else if (num==16'd1753) begin
		AssumePrime = 1;
	end	else if (num==16'd1759) begin
		AssumePrime = 1;
	end	else if (num==16'd1777) begin
		AssumePrime = 1;
	end	else if (num==16'd1783) begin
		AssumePrime = 1;
	end	else if (num==16'd1787) begin
		AssumePrime = 1;
	end	else if (num==16'd1789) begin
		AssumePrime = 1;
	end	else if (num==16'd1801) begin
		AssumePrime = 1;
	end	else if (num==16'd1811) begin
		AssumePrime = 1;
	end	else if (num==16'd1823) begin
		AssumePrime = 1;
	end	else if (num==16'd1831) begin
		AssumePrime = 1;
	end	else if (num==16'd1847) begin
		AssumePrime = 1;
	end	else if (num==16'd1861) begin
		AssumePrime = 1;
	end	else if (num==16'd1867) begin
		AssumePrime = 1;
	end	else if (num==16'd1871) begin
		AssumePrime = 1;
	end	else if (num==16'd1873) begin
		AssumePrime = 1;
	end	else if (num==16'd1877) begin
		AssumePrime = 1;
	end	else if (num==16'd1879) begin
		AssumePrime = 1;
	end	else if (num==16'd1889) begin
		AssumePrime = 1;
	end	else if (num==16'd1901) begin
		AssumePrime = 1;
	end	else if (num==16'd1907) begin
		AssumePrime = 1;
	end	else if (num==16'd1913) begin
		AssumePrime = 1;
	end	else if (num==16'd1931) begin
		AssumePrime = 1;
	end	else if (num==16'd1933) begin
		AssumePrime = 1;
	end	else if (num==16'd1949) begin
		AssumePrime = 1;
	end	else if (num==16'd1951) begin
		AssumePrime = 1;
	end	else if (num==16'd1973) begin
		AssumePrime = 1;
	end	else if (num==16'd1979) begin
		AssumePrime = 1;
	end	else if (num==16'd1987) begin
		AssumePrime = 1;
	end	else if (num==16'd1993) begin
		AssumePrime = 1;
	end	else if (num==16'd1997) begin
		AssumePrime = 1;
	end	else if (num==16'd1999) begin
		AssumePrime = 1;
	end	else if (num==16'd2003) begin
		AssumePrime = 1;
	end	else if (num==16'd2011) begin
		AssumePrime = 1;
	end	else if (num==16'd2017) begin
		AssumePrime = 1;
	end	else if (num==16'd2027) begin
		AssumePrime = 1;
	end	else if (num==16'd2029) begin
		AssumePrime = 1;
	end	else if (num==16'd2039) begin
		AssumePrime = 1;
	end	else if (num==16'd2053) begin
		AssumePrime = 1;
	end	else if (num==16'd2063) begin
		AssumePrime = 1;
	end	else if (num==16'd2069) begin
		AssumePrime = 1;
	end	else if (num==16'd2081) begin
		AssumePrime = 1;
	end	else if (num==16'd2083) begin
		AssumePrime = 1;
	end	else if (num==16'd2087) begin
		AssumePrime = 1;
	end	else if (num==16'd2089) begin
		AssumePrime = 1;
	end	else if (num==16'd2099) begin
		AssumePrime = 1;
	end	else if (num==16'd2111) begin
		AssumePrime = 1;
	end	else if (num==16'd2113) begin
		AssumePrime = 1;
	end	else if (num==16'd2129) begin
		AssumePrime = 1;
	end	else if (num==16'd2131) begin
		AssumePrime = 1;
	end	else if (num==16'd2137) begin
		AssumePrime = 1;
	end	else if (num==16'd2141) begin
		AssumePrime = 1;
	end	else if (num==16'd2143) begin
		AssumePrime = 1;
	end	else if (num==16'd2153) begin
		AssumePrime = 1;
	end	else if (num==16'd2161) begin
		AssumePrime = 1;
	end	else if (num==16'd2179) begin
		AssumePrime = 1;
	end	else if (num==16'd2203) begin
		AssumePrime = 1;
	end	else if (num==16'd2207) begin
		AssumePrime = 1;
	end	else if (num==16'd2213) begin
		AssumePrime = 1;
	end	else if (num==16'd2221) begin
		AssumePrime = 1;
	end	else if (num==16'd2237) begin
		AssumePrime = 1;
	end	else if (num==16'd2239) begin
		AssumePrime = 1;
	end	else if (num==16'd2243) begin
		AssumePrime = 1;
	end	else if (num==16'd2251) begin
		AssumePrime = 1;
	end	else if (num==16'd2267) begin
		AssumePrime = 1;
	end	else if (num==16'd2269) begin
		AssumePrime = 1;
	end	else if (num==16'd2273) begin
		AssumePrime = 1;
	end	else if (num==16'd2281) begin
		AssumePrime = 1;
	end	else if (num==16'd2287) begin
		AssumePrime = 1;
	end	else if (num==16'd2293) begin
		AssumePrime = 1;
	end	else if (num==16'd2297) begin
		AssumePrime = 1;
	end	else if (num==16'd2309) begin
		AssumePrime = 1;
	end	else if (num==16'd2311) begin
		AssumePrime = 1;
	end	else if (num==16'd2333) begin
		AssumePrime = 1;
	end	else if (num==16'd2339) begin
		AssumePrime = 1;
	end	else if (num==16'd2341) begin
		AssumePrime = 1;
	end	else if (num==16'd2347) begin
		AssumePrime = 1;
	end	else if (num==16'd2351) begin
		AssumePrime = 1;
	end	else if (num==16'd2357) begin
		AssumePrime = 1;
	end	else if (num==16'd2371) begin
		AssumePrime = 1;
	end	else if (num==16'd2377) begin
		AssumePrime = 1;
	end	else if (num==16'd2381) begin
		AssumePrime = 1;
	end	else if (num==16'd2383) begin
		AssumePrime = 1;
	end	else if (num==16'd2389) begin
		AssumePrime = 1;
	end	else if (num==16'd2393) begin
		AssumePrime = 1;
	end	else if (num==16'd2399) begin
		AssumePrime = 1;
	end	else if (num==16'd2411) begin
		AssumePrime = 1;
	end	else if (num==16'd2417) begin
		AssumePrime = 1;
	end	else if (num==16'd2423) begin
		AssumePrime = 1;
	end	else if (num==16'd2437) begin
		AssumePrime = 1;
	end	else if (num==16'd2441) begin
		AssumePrime = 1;
	end	else if (num==16'd2447) begin
		AssumePrime = 1;
	end	else if (num==16'd2459) begin
		AssumePrime = 1;
	end	else if (num==16'd2467) begin
		AssumePrime = 1;
	end	else if (num==16'd2473) begin
		AssumePrime = 1;
	end	else if (num==16'd2477) begin
		AssumePrime = 1;
	end	else if (num==16'd2503) begin
		AssumePrime = 1;
	end	else if (num==16'd2521) begin
		AssumePrime = 1;
	end	else if (num==16'd2531) begin
		AssumePrime = 1;
	end	else if (num==16'd2539) begin
		AssumePrime = 1;
	end	else if (num==16'd2543) begin
		AssumePrime = 1;
	end	else if (num==16'd2549) begin
		AssumePrime = 1;
	end	else if (num==16'd2551) begin
		AssumePrime = 1;
	end	else if (num==16'd2557) begin
		AssumePrime = 1;
	end	else if (num==16'd2579) begin
		AssumePrime = 1;
	end	else if (num==16'd2591) begin
		AssumePrime = 1;
	end	else if (num==16'd2593) begin
		AssumePrime = 1;
	end	else if (num==16'd2609) begin
		AssumePrime = 1;
	end	else if (num==16'd2617) begin
		AssumePrime = 1;
	end	else if (num==16'd2621) begin
		AssumePrime = 1;
	end	else if (num==16'd2633) begin
		AssumePrime = 1;
	end	else if (num==16'd2647) begin
		AssumePrime = 1;
	end	else if (num==16'd2657) begin
		AssumePrime = 1;
	end	else if (num==16'd2659) begin
		AssumePrime = 1;
	end	else if (num==16'd2663) begin
		AssumePrime = 1;
	end	else if (num==16'd2671) begin
		AssumePrime = 1;
	end	else if (num==16'd2677) begin
		AssumePrime = 1;
	end	else if (num==16'd2683) begin
		AssumePrime = 1;
	end	else if (num==16'd2687) begin
		AssumePrime = 1;
	end	else if (num==16'd2689) begin
		AssumePrime = 1;
	end	else if (num==16'd2693) begin
		AssumePrime = 1;
	end	else if (num==16'd2699) begin
		AssumePrime = 1;
	end	else if (num==16'd2707) begin
		AssumePrime = 1;
	end	else if (num==16'd2711) begin
		AssumePrime = 1;
	end	else if (num==16'd2713) begin
		AssumePrime = 1;
	end	else if (num==16'd2719) begin
		AssumePrime = 1;
	end	else if (num==16'd2729) begin
		AssumePrime = 1;
	end	else if (num==16'd2731) begin
		AssumePrime = 1;
	end	else if (num==16'd2741) begin
		AssumePrime = 1;
	end	else if (num==16'd2749) begin
		AssumePrime = 1;
	end	else if (num==16'd2753) begin
		AssumePrime = 1;
	end	else if (num==16'd2767) begin
		AssumePrime = 1;
	end	else if (num==16'd2777) begin
		AssumePrime = 1;
	end	else if (num==16'd2789) begin
		AssumePrime = 1;
	end	else if (num==16'd2791) begin
		AssumePrime = 1;
	end	else if (num==16'd2797) begin
		AssumePrime = 1;
	end	else if (num==16'd2801) begin
		AssumePrime = 1;
	end	else if (num==16'd2803) begin
		AssumePrime = 1;
	end	else if (num==16'd2819) begin
		AssumePrime = 1;
	end	else if (num==16'd2833) begin
		AssumePrime = 1;
	end	else if (num==16'd2837) begin
		AssumePrime = 1;
	end	else if (num==16'd2843) begin
		AssumePrime = 1;
	end	else if (num==16'd2851) begin
		AssumePrime = 1;
	end	else if (num==16'd2857) begin
		AssumePrime = 1;
	end	else if (num==16'd2861) begin
		AssumePrime = 1;
	end	else if (num==16'd2879) begin
		AssumePrime = 1;
	end	else if (num==16'd2887) begin
		AssumePrime = 1;
	end	else if (num==16'd2897) begin
		AssumePrime = 1;
	end	else if (num==16'd2903) begin
		AssumePrime = 1;
	end	else if (num==16'd2909) begin
		AssumePrime = 1;
	end	else if (num==16'd2917) begin
		AssumePrime = 1;
	end	else if (num==16'd2927) begin
		AssumePrime = 1;
	end	else if (num==16'd2939) begin
		AssumePrime = 1;
	end	else if (num==16'd2953) begin
		AssumePrime = 1;
	end	else if (num==16'd2957) begin
		AssumePrime = 1;
	end	else if (num==16'd2963) begin
		AssumePrime = 1;
	end	else if (num==16'd2969) begin
		AssumePrime = 1;
	end	else if (num==16'd2971) begin
		AssumePrime = 1;
	end	else if (num==16'd2999) begin
		AssumePrime = 1;
	end	else if (num==16'd3001) begin
		AssumePrime = 1;
	end	else if (num==16'd3011) begin
		AssumePrime = 1;
	end	else if (num==16'd3019) begin
		AssumePrime = 1;
	end	else if (num==16'd3023) begin
		AssumePrime = 1;
	end	else if (num==16'd3037) begin
		AssumePrime = 1;
	end	else if (num==16'd3041) begin
		AssumePrime = 1;
	end	else if (num==16'd3049) begin
		AssumePrime = 1;
	end	else if (num==16'd3061) begin
		AssumePrime = 1;
	end	else if (num==16'd3067) begin
		AssumePrime = 1;
	end	else if (num==16'd3079) begin
		AssumePrime = 1;
	end	else if (num==16'd3083) begin
		AssumePrime = 1;
	end	else if (num==16'd3089) begin
		AssumePrime = 1;
	end	else if (num==16'd3109) begin
		AssumePrime = 1;
	end	else if (num==16'd3119) begin
		AssumePrime = 1;
	end	else if (num==16'd3121) begin
		AssumePrime = 1;
	end	else if (num==16'd3137) begin
		AssumePrime = 1;
	end	else if (num==16'd3163) begin
		AssumePrime = 1;
	end	else if (num==16'd3167) begin
		AssumePrime = 1;
	end	else if (num==16'd3169) begin
		AssumePrime = 1;
	end	else if (num==16'd3181) begin
		AssumePrime = 1;
	end	else if (num==16'd3187) begin
		AssumePrime = 1;
	end	else if (num==16'd3191) begin
		AssumePrime = 1;
	end	else if (num==16'd3203) begin
		AssumePrime = 1;
	end	else if (num==16'd3209) begin
		AssumePrime = 1;
	end	else if (num==16'd3217) begin
		AssumePrime = 1;
	end	else if (num==16'd3221) begin
		AssumePrime = 1;
	end	else if (num==16'd3229) begin
		AssumePrime = 1;
	end	else if (num==16'd3251) begin
		AssumePrime = 1;
	end	else if (num==16'd3253) begin
		AssumePrime = 1;
	end	else if (num==16'd3257) begin
		AssumePrime = 1;
	end	else if (num==16'd3259) begin
		AssumePrime = 1;
	end	else if (num==16'd3271) begin
		AssumePrime = 1;
	end	else if (num==16'd3299) begin
		AssumePrime = 1;
	end	else if (num==16'd3301) begin
		AssumePrime = 1;
	end	else if (num==16'd3307) begin
		AssumePrime = 1;
	end	else if (num==16'd3313) begin
		AssumePrime = 1;
	end	else if (num==16'd3319) begin
		AssumePrime = 1;
	end	else if (num==16'd3323) begin
		AssumePrime = 1;
	end	else if (num==16'd3329) begin
		AssumePrime = 1;
	end	else if (num==16'd3331) begin
		AssumePrime = 1;
	end	else if (num==16'd3343) begin
		AssumePrime = 1;
	end	else if (num==16'd3347) begin
		AssumePrime = 1;
	end	else if (num==16'd3359) begin
		AssumePrime = 1;
	end	else if (num==16'd3361) begin
		AssumePrime = 1;
	end	else if (num==16'd3371) begin
		AssumePrime = 1;
	end	else if (num==16'd3373) begin
		AssumePrime = 1;
	end	else if (num==16'd3389) begin
		AssumePrime = 1;
	end	else if (num==16'd3391) begin
		AssumePrime = 1;
	end	else if (num==16'd3407) begin
		AssumePrime = 1;
	end	else if (num==16'd3413) begin
		AssumePrime = 1;
	end	else if (num==16'd3433) begin
		AssumePrime = 1;
	end	else if (num==16'd3449) begin
		AssumePrime = 1;
	end	else if (num==16'd3457) begin
		AssumePrime = 1;
	end	else if (num==16'd3461) begin
		AssumePrime = 1;
	end	else if (num==16'd3463) begin
		AssumePrime = 1;
	end	else if (num==16'd3467) begin
		AssumePrime = 1;
	end	else if (num==16'd3469) begin
		AssumePrime = 1;
	end	else if (num==16'd3491) begin
		AssumePrime = 1;
	end	else if (num==16'd3499) begin
		AssumePrime = 1;
	end	else if (num==16'd3511) begin
		AssumePrime = 1;
	end	else if (num==16'd3517) begin
		AssumePrime = 1;
	end	else if (num==16'd3527) begin
		AssumePrime = 1;
	end	else if (num==16'd3529) begin
		AssumePrime = 1;
	end	else if (num==16'd3533) begin
		AssumePrime = 1;
	end	else if (num==16'd3539) begin
		AssumePrime = 1;
	end	else if (num==16'd3541) begin
		AssumePrime = 1;
	end	else if (num==16'd3547) begin
		AssumePrime = 1;
	end	else if (num==16'd3557) begin
		AssumePrime = 1;
	end	else if (num==16'd3559) begin
		AssumePrime = 1;
	end	else if (num==16'd3571) begin
		AssumePrime = 1;
	end	else if (num==16'd3581) begin
		AssumePrime = 1;
	end	else if (num==16'd3583) begin
		AssumePrime = 1;
	end	else if (num==16'd3593) begin
		AssumePrime = 1;
	end	else if (num==16'd3607) begin
		AssumePrime = 1;
	end	else if (num==16'd3613) begin
		AssumePrime = 1;
	end	else if (num==16'd3617) begin
		AssumePrime = 1;
	end	else if (num==16'd3623) begin
		AssumePrime = 1;
	end	else if (num==16'd3631) begin
		AssumePrime = 1;
	end	else if (num==16'd3637) begin
		AssumePrime = 1;
	end	else if (num==16'd3643) begin
		AssumePrime = 1;
	end	else if (num==16'd3659) begin
		AssumePrime = 1;
	end	else if (num==16'd3671) begin
		AssumePrime = 1;
	end	else if (num==16'd3673) begin
		AssumePrime = 1;
	end	else if (num==16'd3677) begin
		AssumePrime = 1;
	end	else if (num==16'd3691) begin
		AssumePrime = 1;
	end	else if (num==16'd3697) begin
		AssumePrime = 1;
	end	else if (num==16'd3701) begin
		AssumePrime = 1;
	end	else if (num==16'd3709) begin
		AssumePrime = 1;
	end	else if (num==16'd3719) begin
		AssumePrime = 1;
	end	else if (num==16'd3727) begin
		AssumePrime = 1;
	end	else if (num==16'd3733) begin
		AssumePrime = 1;
	end	else if (num==16'd3739) begin
		AssumePrime = 1;
	end	else if (num==16'd3761) begin
		AssumePrime = 1;
	end	else if (num==16'd3767) begin
		AssumePrime = 1;
	end	else if (num==16'd3769) begin
		AssumePrime = 1;
	end	else if (num==16'd3779) begin
		AssumePrime = 1;
	end	else if (num==16'd3793) begin
		AssumePrime = 1;
	end	else if (num==16'd3797) begin
		AssumePrime = 1;
	end	else if (num==16'd3803) begin
		AssumePrime = 1;
	end	else if (num==16'd3821) begin
		AssumePrime = 1;
	end	else if (num==16'd3823) begin
		AssumePrime = 1;
	end	else if (num==16'd3833) begin
		AssumePrime = 1;
	end	else if (num==16'd3847) begin
		AssumePrime = 1;
	end	else if (num==16'd3851) begin
		AssumePrime = 1;
	end	else if (num==16'd3853) begin
		AssumePrime = 1;
	end	else if (num==16'd3863) begin
		AssumePrime = 1;
	end	else if (num==16'd3877) begin
		AssumePrime = 1;
	end	else if (num==16'd3881) begin
		AssumePrime = 1;
	end	else if (num==16'd3889) begin
		AssumePrime = 1;
	end	else if (num==16'd3907) begin
		AssumePrime = 1;
	end	else if (num==16'd3911) begin
		AssumePrime = 1;
	end	else if (num==16'd3917) begin
		AssumePrime = 1;
	end	else if (num==16'd3919) begin
		AssumePrime = 1;
	end	else if (num==16'd3923) begin
		AssumePrime = 1;
	end	else if (num==16'd3929) begin
		AssumePrime = 1;
	end	else if (num==16'd3931) begin
		AssumePrime = 1;
	end	else if (num==16'd3943) begin
		AssumePrime = 1;
	end	else if (num==16'd3947) begin
		AssumePrime = 1;
	end	else if (num==16'd3967) begin
		AssumePrime = 1;
	end	else if (num==16'd3989) begin
		AssumePrime = 1;
	end	else if (num==16'd4001) begin
		AssumePrime = 1;
	end	else if (num==16'd4003) begin
		AssumePrime = 1;
	end	else if (num==16'd4007) begin
		AssumePrime = 1;
	end	else if (num==16'd4013) begin
		AssumePrime = 1;
	end	else if (num==16'd4019) begin
		AssumePrime = 1;
	end	else if (num==16'd4021) begin
		AssumePrime = 1;
	end	else if (num==16'd4027) begin
		AssumePrime = 1;
	end	else if (num==16'd4049) begin
		AssumePrime = 1;
	end	else if (num==16'd4051) begin
		AssumePrime = 1;
	end	else if (num==16'd4057) begin
		AssumePrime = 1;
	end	else if (num==16'd4073) begin
		AssumePrime = 1;
	end	else if (num==16'd4079) begin
		AssumePrime = 1;
	end	else if (num==16'd4091) begin
		AssumePrime = 1;
	end	else if (num==16'd4093) begin
		AssumePrime = 1;
	end	else if (num==16'd4099) begin
		AssumePrime = 1;
	end	else if (num==16'd4111) begin
		AssumePrime = 1;
	end	else if (num==16'd4127) begin
		AssumePrime = 1;
	end	else if (num==16'd4129) begin
		AssumePrime = 1;
	end	else if (num==16'd4133) begin
		AssumePrime = 1;
	end	else if (num==16'd4139) begin
		AssumePrime = 1;
	end	else if (num==16'd4153) begin
		AssumePrime = 1;
	end	else if (num==16'd4157) begin
		AssumePrime = 1;
	end	else if (num==16'd4159) begin
		AssumePrime = 1;
	end	else if (num==16'd4177) begin
		AssumePrime = 1;
	end	else if (num==16'd4201) begin
		AssumePrime = 1;
	end	else if (num==16'd4211) begin
		AssumePrime = 1;
	end	else if (num==16'd4217) begin
		AssumePrime = 1;
	end	else if (num==16'd4219) begin
		AssumePrime = 1;
	end	else if (num==16'd4229) begin
		AssumePrime = 1;
	end	else if (num==16'd4231) begin
		AssumePrime = 1;
	end	else if (num==16'd4241) begin
		AssumePrime = 1;
	end	else if (num==16'd4243) begin
		AssumePrime = 1;
	end	else if (num==16'd4253) begin
		AssumePrime = 1;
	end	else if (num==16'd4259) begin
		AssumePrime = 1;
	end	else if (num==16'd4261) begin
		AssumePrime = 1;
	end	else if (num==16'd4271) begin
		AssumePrime = 1;
	end	else if (num==16'd4273) begin
		AssumePrime = 1;
	end	else if (num==16'd4283) begin
		AssumePrime = 1;
	end	else if (num==16'd4289) begin
		AssumePrime = 1;
	end	else if (num==16'd4297) begin
		AssumePrime = 1;
	end	else if (num==16'd4327) begin
		AssumePrime = 1;
	end	else if (num==16'd4337) begin
		AssumePrime = 1;
	end	else if (num==16'd4339) begin
		AssumePrime = 1;
	end	else if (num==16'd4349) begin
		AssumePrime = 1;
	end	else if (num==16'd4357) begin
		AssumePrime = 1;
	end	else if (num==16'd4363) begin
		AssumePrime = 1;
	end	else if (num==16'd4373) begin
		AssumePrime = 1;
	end	else if (num==16'd4391) begin
		AssumePrime = 1;
	end	else if (num==16'd4397) begin
		AssumePrime = 1;
	end	else if (num==16'd4409) begin
		AssumePrime = 1;
	end	else if (num==16'd4421) begin
		AssumePrime = 1;
	end	else if (num==16'd4423) begin
		AssumePrime = 1;
	end	else if (num==16'd4441) begin
		AssumePrime = 1;
	end	else if (num==16'd4447) begin
		AssumePrime = 1;
	end	else if (num==16'd4451) begin
		AssumePrime = 1;
	end	else if (num==16'd4457) begin
		AssumePrime = 1;
	end	else if (num==16'd4463) begin
		AssumePrime = 1;
	end	else if (num==16'd4481) begin
		AssumePrime = 1;
	end	else if (num==16'd4483) begin
		AssumePrime = 1;
	end	else if (num==16'd4493) begin
		AssumePrime = 1;
	end	else if (num==16'd4507) begin
		AssumePrime = 1;
	end	else if (num==16'd4513) begin
		AssumePrime = 1;
	end	else if (num==16'd4517) begin
		AssumePrime = 1;
	end	else if (num==16'd4519) begin
		AssumePrime = 1;
	end	else if (num==16'd4523) begin
		AssumePrime = 1;
	end	else if (num==16'd4547) begin
		AssumePrime = 1;
	end	else if (num==16'd4549) begin
		AssumePrime = 1;
	end	else if (num==16'd4561) begin
		AssumePrime = 1;
	end	else if (num==16'd4567) begin
		AssumePrime = 1;
	end	else if (num==16'd4583) begin
		AssumePrime = 1;
	end	else if (num==16'd4591) begin
		AssumePrime = 1;
	end	else if (num==16'd4597) begin
		AssumePrime = 1;
	end	else if (num==16'd4603) begin
		AssumePrime = 1;
	end	else if (num==16'd4621) begin
		AssumePrime = 1;
	end	else if (num==16'd4637) begin
		AssumePrime = 1;
	end	else if (num==16'd4639) begin
		AssumePrime = 1;
	end	else if (num==16'd4643) begin
		AssumePrime = 1;
	end	else if (num==16'd4649) begin
		AssumePrime = 1;
	end	else if (num==16'd4651) begin
		AssumePrime = 1;
	end	else if (num==16'd4657) begin
		AssumePrime = 1;
	end	else if (num==16'd4663) begin
		AssumePrime = 1;
	end	else if (num==16'd4673) begin
		AssumePrime = 1;
	end	else if (num==16'd4679) begin
		AssumePrime = 1;
	end	else if (num==16'd4691) begin
		AssumePrime = 1;
	end	else if (num==16'd4703) begin
		AssumePrime = 1;
	end	else if (num==16'd4721) begin
		AssumePrime = 1;
	end	else if (num==16'd4723) begin
		AssumePrime = 1;
	end	else if (num==16'd4729) begin
		AssumePrime = 1;
	end	else if (num==16'd4733) begin
		AssumePrime = 1;
	end	else if (num==16'd4751) begin
		AssumePrime = 1;
	end	else if (num==16'd4759) begin
		AssumePrime = 1;
	end	else if (num==16'd4783) begin
		AssumePrime = 1;
	end	else if (num==16'd4787) begin
		AssumePrime = 1;
	end	else if (num==16'd4789) begin
		AssumePrime = 1;
	end	else if (num==16'd4793) begin
		AssumePrime = 1;
	end	else if (num==16'd4799) begin
		AssumePrime = 1;
	end	else if (num==16'd4801) begin
		AssumePrime = 1;
	end	else if (num==16'd4813) begin
		AssumePrime = 1;
	end	else if (num==16'd4817) begin
		AssumePrime = 1;
	end	else if (num==16'd4831) begin
		AssumePrime = 1;
	end	else if (num==16'd4861) begin
		AssumePrime = 1;
	end	else if (num==16'd4871) begin
		AssumePrime = 1;
	end	else if (num==16'd4877) begin
		AssumePrime = 1;
	end	else if (num==16'd4889) begin
		AssumePrime = 1;
	end	else if (num==16'd4903) begin
		AssumePrime = 1;
	end	else if (num==16'd4909) begin
		AssumePrime = 1;
	end	else if (num==16'd4919) begin
		AssumePrime = 1;
	end	else if (num==16'd4931) begin
		AssumePrime = 1;
	end	else if (num==16'd4933) begin
		AssumePrime = 1;
	end	else if (num==16'd4937) begin
		AssumePrime = 1;
	end	else if (num==16'd4943) begin
		AssumePrime = 1;
	end	else if (num==16'd4951) begin
		AssumePrime = 1;
	end	else if (num==16'd4957) begin
		AssumePrime = 1;
	end	else if (num==16'd4967) begin
		AssumePrime = 1;
	end	else if (num==16'd4969) begin
		AssumePrime = 1;
	end	else if (num==16'd4973) begin
		AssumePrime = 1;
	end	else if (num==16'd4987) begin
		AssumePrime = 1;
	end	else if (num==16'd4993) begin
		AssumePrime = 1;
	end	else if (num==16'd4999) begin
		AssumePrime = 1;
	end	else if (num==16'd5003) begin
		AssumePrime = 1;
	end	else if (num==16'd5009) begin
		AssumePrime = 1;
	end	else if (num==16'd5011) begin
		AssumePrime = 1;
	end	else if (num==16'd5021) begin
		AssumePrime = 1;
	end	else if (num==16'd5023) begin
		AssumePrime = 1;
	end	else if (num==16'd5039) begin
		AssumePrime = 1;
	end	else if (num==16'd5051) begin
		AssumePrime = 1;
	end	else if (num==16'd5059) begin
		AssumePrime = 1;
	end	else if (num==16'd5077) begin
		AssumePrime = 1;
	end	else if (num==16'd5081) begin
		AssumePrime = 1;
	end	else if (num==16'd5087) begin
		AssumePrime = 1;
	end	else if (num==16'd5099) begin
		AssumePrime = 1;
	end	else if (num==16'd5101) begin
		AssumePrime = 1;
	end	else if (num==16'd5107) begin
		AssumePrime = 1;
	end	else if (num==16'd5113) begin
		AssumePrime = 1;
	end	else if (num==16'd5119) begin
		AssumePrime = 1;
	end	else if (num==16'd5147) begin
		AssumePrime = 1;
	end	else if (num==16'd5153) begin
		AssumePrime = 1;
	end	else if (num==16'd5167) begin
		AssumePrime = 1;
	end	else if (num==16'd5171) begin
		AssumePrime = 1;
	end	else if (num==16'd5179) begin
		AssumePrime = 1;
	end	else if (num==16'd5189) begin
		AssumePrime = 1;
	end	else if (num==16'd5197) begin
		AssumePrime = 1;
	end	else if (num==16'd5209) begin
		AssumePrime = 1;
	end	else if (num==16'd5227) begin
		AssumePrime = 1;
	end	else if (num==16'd5231) begin
		AssumePrime = 1;
	end	else if (num==16'd5233) begin
		AssumePrime = 1;
	end	else if (num==16'd5237) begin
		AssumePrime = 1;
	end	else if (num==16'd5261) begin
		AssumePrime = 1;
	end	else if (num==16'd5273) begin
		AssumePrime = 1;
	end	else if (num==16'd5279) begin
		AssumePrime = 1;
	end	else if (num==16'd5281) begin
		AssumePrime = 1;
	end	else if (num==16'd5297) begin
		AssumePrime = 1;
	end	else if (num==16'd5303) begin
		AssumePrime = 1;
	end	else if (num==16'd5309) begin
		AssumePrime = 1;
	end	else if (num==16'd5323) begin
		AssumePrime = 1;
	end	else if (num==16'd5333) begin
		AssumePrime = 1;
	end	else if (num==16'd5347) begin
		AssumePrime = 1;
	end	else if (num==16'd5351) begin
		AssumePrime = 1;
	end	else if (num==16'd5381) begin
		AssumePrime = 1;
	end	else if (num==16'd5387) begin
		AssumePrime = 1;
	end	else if (num==16'd5393) begin
		AssumePrime = 1;
	end	else if (num==16'd5399) begin
		AssumePrime = 1;
	end	else if (num==16'd5407) begin
		AssumePrime = 1;
	end	else if (num==16'd5413) begin
		AssumePrime = 1;
	end	else if (num==16'd5417) begin
		AssumePrime = 1;
	end	else if (num==16'd5419) begin
		AssumePrime = 1;
	end	else if (num==16'd5431) begin
		AssumePrime = 1;
	end	else if (num==16'd5437) begin
		AssumePrime = 1;
	end	else if (num==16'd5441) begin
		AssumePrime = 1;
	end	else if (num==16'd5443) begin
		AssumePrime = 1;
	end	else if (num==16'd5449) begin
		AssumePrime = 1;
	end	else if (num==16'd5471) begin
		AssumePrime = 1;
	end	else if (num==16'd5477) begin
		AssumePrime = 1;
	end	else if (num==16'd5479) begin
		AssumePrime = 1;
	end	else if (num==16'd5483) begin
		AssumePrime = 1;
	end	else if (num==16'd5501) begin
		AssumePrime = 1;
	end	else if (num==16'd5503) begin
		AssumePrime = 1;
	end	else if (num==16'd5507) begin
		AssumePrime = 1;
	end	else if (num==16'd5519) begin
		AssumePrime = 1;
	end	else if (num==16'd5521) begin
		AssumePrime = 1;
	end	else if (num==16'd5527) begin
		AssumePrime = 1;
	end	else if (num==16'd5531) begin
		AssumePrime = 1;
	end	else if (num==16'd5557) begin
		AssumePrime = 1;
	end	else if (num==16'd5563) begin
		AssumePrime = 1;
	end	else if (num==16'd5569) begin
		AssumePrime = 1;
	end	else if (num==16'd5573) begin
		AssumePrime = 1;
	end	else if (num==16'd5581) begin
		AssumePrime = 1;
	end	else if (num==16'd5591) begin
		AssumePrime = 1;
	end	else if (num==16'd5623) begin
		AssumePrime = 1;
	end	else if (num==16'd5639) begin
		AssumePrime = 1;
	end	else if (num==16'd5641) begin
		AssumePrime = 1;
	end	else if (num==16'd5647) begin
		AssumePrime = 1;
	end	else if (num==16'd5651) begin
		AssumePrime = 1;
	end	else if (num==16'd5653) begin
		AssumePrime = 1;
	end	else if (num==16'd5657) begin
		AssumePrime = 1;
	end	else if (num==16'd5659) begin
		AssumePrime = 1;
	end	else if (num==16'd5669) begin
		AssumePrime = 1;
	end	else if (num==16'd5683) begin
		AssumePrime = 1;
	end	else if (num==16'd5689) begin
		AssumePrime = 1;
	end	else if (num==16'd5693) begin
		AssumePrime = 1;
	end	else if (num==16'd5701) begin
		AssumePrime = 1;
	end	else if (num==16'd5711) begin
		AssumePrime = 1;
	end	else if (num==16'd5717) begin
		AssumePrime = 1;
	end	else if (num==16'd5737) begin
		AssumePrime = 1;
	end	else if (num==16'd5741) begin
		AssumePrime = 1;
	end	else if (num==16'd5743) begin
		AssumePrime = 1;
	end	else if (num==16'd5749) begin
		AssumePrime = 1;
	end	else if (num==16'd5779) begin
		AssumePrime = 1;
	end	else if (num==16'd5783) begin
		AssumePrime = 1;
	end	else if (num==16'd5791) begin
		AssumePrime = 1;
	end	else if (num==16'd5801) begin
		AssumePrime = 1;
	end	else if (num==16'd5807) begin
		AssumePrime = 1;
	end	else if (num==16'd5813) begin
		AssumePrime = 1;
	end	else if (num==16'd5821) begin
		AssumePrime = 1;
	end	else if (num==16'd5827) begin
		AssumePrime = 1;
	end	else if (num==16'd5839) begin
		AssumePrime = 1;
	end	else if (num==16'd5843) begin
		AssumePrime = 1;
	end	else if (num==16'd5849) begin
		AssumePrime = 1;
	end	else if (num==16'd5851) begin
		AssumePrime = 1;
	end	else if (num==16'd5857) begin
		AssumePrime = 1;
	end	else if (num==16'd5861) begin
		AssumePrime = 1;
	end	else if (num==16'd5867) begin
		AssumePrime = 1;
	end	else if (num==16'd5869) begin
		AssumePrime = 1;
	end	else if (num==16'd5879) begin
		AssumePrime = 1;
	end	else if (num==16'd5881) begin
		AssumePrime = 1;
	end	else if (num==16'd5897) begin
		AssumePrime = 1;
	end	else if (num==16'd5903) begin
		AssumePrime = 1;
	end	else if (num==16'd5923) begin
		AssumePrime = 1;
	end	else if (num==16'd5927) begin
		AssumePrime = 1;
	end	else if (num==16'd5939) begin
		AssumePrime = 1;
	end	else if (num==16'd5953) begin
		AssumePrime = 1;
	end	else if (num==16'd5981) begin
		AssumePrime = 1;
	end	else if (num==16'd5987) begin
		AssumePrime = 1;
	end	else if (num==16'd6007) begin
		AssumePrime = 1;
	end	else if (num==16'd6011) begin
		AssumePrime = 1;
	end	else if (num==16'd6029) begin
		AssumePrime = 1;
	end	else if (num==16'd6037) begin
		AssumePrime = 1;
	end	else if (num==16'd6043) begin
		AssumePrime = 1;
	end	else if (num==16'd6047) begin
		AssumePrime = 1;
	end	else if (num==16'd6053) begin
		AssumePrime = 1;
	end	else if (num==16'd6067) begin
		AssumePrime = 1;
	end	else if (num==16'd6073) begin
		AssumePrime = 1;
	end	else if (num==16'd6079) begin
		AssumePrime = 1;
	end	else if (num==16'd6089) begin
		AssumePrime = 1;
	end	else if (num==16'd6091) begin
		AssumePrime = 1;
	end	else if (num==16'd6101) begin
		AssumePrime = 1;
	end	else if (num==16'd6113) begin
		AssumePrime = 1;
	end	else if (num==16'd6121) begin
		AssumePrime = 1;
	end	else if (num==16'd6131) begin
		AssumePrime = 1;
	end	else if (num==16'd6133) begin
		AssumePrime = 1;
	end	else if (num==16'd6143) begin
		AssumePrime = 1;
	end	else if (num==16'd6151) begin
		AssumePrime = 1;
	end	else if (num==16'd6163) begin
		AssumePrime = 1;
	end	else if (num==16'd6173) begin
		AssumePrime = 1;
	end	else if (num==16'd6197) begin
		AssumePrime = 1;
	end	else if (num==16'd6199) begin
		AssumePrime = 1;
	end	else if (num==16'd6203) begin
		AssumePrime = 1;
	end	else if (num==16'd6211) begin
		AssumePrime = 1;
	end	else if (num==16'd6217) begin
		AssumePrime = 1;
	end	else if (num==16'd6221) begin
		AssumePrime = 1;
	end	else if (num==16'd6229) begin
		AssumePrime = 1;
	end	else if (num==16'd6247) begin
		AssumePrime = 1;
	end	else if (num==16'd6257) begin
		AssumePrime = 1;
	end	else if (num==16'd6263) begin
		AssumePrime = 1;
	end	else if (num==16'd6269) begin
		AssumePrime = 1;
	end	else if (num==16'd6271) begin
		AssumePrime = 1;
	end	else if (num==16'd6277) begin
		AssumePrime = 1;
	end	else if (num==16'd6287) begin
		AssumePrime = 1;
	end	else if (num==16'd6299) begin
		AssumePrime = 1;
	end	else if (num==16'd6301) begin
		AssumePrime = 1;
	end	else if (num==16'd6311) begin
		AssumePrime = 1;
	end	else if (num==16'd6317) begin
		AssumePrime = 1;
	end	else if (num==16'd6323) begin
		AssumePrime = 1;
	end	else if (num==16'd6329) begin
		AssumePrime = 1;
	end	else if (num==16'd6337) begin
		AssumePrime = 1;
	end	else if (num==16'd6343) begin
		AssumePrime = 1;
	end	else if (num==16'd6353) begin
		AssumePrime = 1;
	end	else if (num==16'd6359) begin
		AssumePrime = 1;
	end	else if (num==16'd6361) begin
		AssumePrime = 1;
	end	else if (num==16'd6367) begin
		AssumePrime = 1;
	end	else if (num==16'd6373) begin
		AssumePrime = 1;
	end	else if (num==16'd6379) begin
		AssumePrime = 1;
	end	else if (num==16'd6389) begin
		AssumePrime = 1;
	end	else if (num==16'd6397) begin
		AssumePrime = 1;
	end	else if (num==16'd6421) begin
		AssumePrime = 1;
	end	else if (num==16'd6427) begin
		AssumePrime = 1;
	end	else if (num==16'd6449) begin
		AssumePrime = 1;
	end	else if (num==16'd6451) begin
		AssumePrime = 1;
	end	else if (num==16'd6469) begin
		AssumePrime = 1;
	end	else if (num==16'd6473) begin
		AssumePrime = 1;
	end	else if (num==16'd6481) begin
		AssumePrime = 1;
	end	else if (num==16'd6491) begin
		AssumePrime = 1;
	end	else if (num==16'd6521) begin
		AssumePrime = 1;
	end	else if (num==16'd6529) begin
		AssumePrime = 1;
	end	else if (num==16'd6547) begin
		AssumePrime = 1;
	end	else if (num==16'd6551) begin
		AssumePrime = 1;
	end	else if (num==16'd6553) begin
		AssumePrime = 1;
	end	else if (num==16'd6563) begin
		AssumePrime = 1;
	end	else if (num==16'd6569) begin
		AssumePrime = 1;
	end	else if (num==16'd6571) begin
		AssumePrime = 1;
	end	else if (num==16'd6577) begin
		AssumePrime = 1;
	end	else if (num==16'd6581) begin
		AssumePrime = 1;
	end	else if (num==16'd6599) begin
		AssumePrime = 1;
	end	else if (num==16'd6607) begin
		AssumePrime = 1;
	end	else if (num==16'd6619) begin
		AssumePrime = 1;
	end	else if (num==16'd6637) begin
		AssumePrime = 1;
	end	else if (num==16'd6653) begin
		AssumePrime = 1;
	end	else if (num==16'd6659) begin
		AssumePrime = 1;
	end	else if (num==16'd6661) begin
		AssumePrime = 1;
	end	else if (num==16'd6673) begin
		AssumePrime = 1;
	end	else if (num==16'd6679) begin
		AssumePrime = 1;
	end	else if (num==16'd6689) begin
		AssumePrime = 1;
	end	else if (num==16'd6691) begin
		AssumePrime = 1;
	end	else if (num==16'd6701) begin
		AssumePrime = 1;
	end	else if (num==16'd6703) begin
		AssumePrime = 1;
	end	else if (num==16'd6709) begin
		AssumePrime = 1;
	end	else if (num==16'd6719) begin
		AssumePrime = 1;
	end	else if (num==16'd6733) begin
		AssumePrime = 1;
	end	else if (num==16'd6737) begin
		AssumePrime = 1;
	end	else if (num==16'd6761) begin
		AssumePrime = 1;
	end	else if (num==16'd6763) begin
		AssumePrime = 1;
	end	else if (num==16'd6779) begin
		AssumePrime = 1;
	end	else if (num==16'd6781) begin
		AssumePrime = 1;
	end	else if (num==16'd6791) begin
		AssumePrime = 1;
	end	else if (num==16'd6793) begin
		AssumePrime = 1;
	end	else if (num==16'd6803) begin
		AssumePrime = 1;
	end	else if (num==16'd6823) begin
		AssumePrime = 1;
	end	else if (num==16'd6827) begin
		AssumePrime = 1;
	end	else if (num==16'd6829) begin
		AssumePrime = 1;
	end	else if (num==16'd6833) begin
		AssumePrime = 1;
	end	else if (num==16'd6841) begin
		AssumePrime = 1;
	end	else if (num==16'd6857) begin
		AssumePrime = 1;
	end	else if (num==16'd6863) begin
		AssumePrime = 1;
	end	else if (num==16'd6869) begin
		AssumePrime = 1;
	end	else if (num==16'd6871) begin
		AssumePrime = 1;
	end	else if (num==16'd6883) begin
		AssumePrime = 1;
	end	else if (num==16'd6899) begin
		AssumePrime = 1;
	end	else if (num==16'd6907) begin
		AssumePrime = 1;
	end	else if (num==16'd6911) begin
		AssumePrime = 1;
	end	else if (num==16'd6917) begin
		AssumePrime = 1;
	end	else if (num==16'd6947) begin
		AssumePrime = 1;
	end	else if (num==16'd6949) begin
		AssumePrime = 1;
	end	else if (num==16'd6959) begin
		AssumePrime = 1;
	end	else if (num==16'd6961) begin
		AssumePrime = 1;
	end	else if (num==16'd6967) begin
		AssumePrime = 1;
	end	else if (num==16'd6971) begin
		AssumePrime = 1;
	end	else if (num==16'd6977) begin
		AssumePrime = 1;
	end	else if (num==16'd6983) begin
		AssumePrime = 1;
	end	else if (num==16'd6991) begin
		AssumePrime = 1;
	end	else if (num==16'd6997) begin
		AssumePrime = 1;
	end	else if (num==16'd7001) begin
		AssumePrime = 1;
	end	else if (num==16'd7013) begin
		AssumePrime = 1;
	end	else if (num==16'd7019) begin
		AssumePrime = 1;
	end	else if (num==16'd7027) begin
		AssumePrime = 1;
	end	else if (num==16'd7039) begin
		AssumePrime = 1;
	end	else if (num==16'd7043) begin
		AssumePrime = 1;
	end	else if (num==16'd7057) begin
		AssumePrime = 1;
	end	else if (num==16'd7069) begin
		AssumePrime = 1;
	end	else if (num==16'd7079) begin
		AssumePrime = 1;
	end	else if (num==16'd7103) begin
		AssumePrime = 1;
	end	else if (num==16'd7109) begin
		AssumePrime = 1;
	end	else if (num==16'd7121) begin
		AssumePrime = 1;
	end	else if (num==16'd7127) begin
		AssumePrime = 1;
	end	else if (num==16'd7129) begin
		AssumePrime = 1;
	end	else if (num==16'd7151) begin
		AssumePrime = 1;
	end	else if (num==16'd7159) begin
		AssumePrime = 1;
	end	else if (num==16'd7177) begin
		AssumePrime = 1;
	end	else if (num==16'd7187) begin
		AssumePrime = 1;
	end	else if (num==16'd7193) begin
		AssumePrime = 1;
	end	else if (num==16'd7207) begin
		AssumePrime = 1;
	end	else if (num==16'd7211) begin
		AssumePrime = 1;
	end	else if (num==16'd7213) begin
		AssumePrime = 1;
	end	else if (num==16'd7219) begin
		AssumePrime = 1;
	end	else if (num==16'd7229) begin
		AssumePrime = 1;
	end	else if (num==16'd7237) begin
		AssumePrime = 1;
	end	else if (num==16'd7243) begin
		AssumePrime = 1;
	end	else if (num==16'd7247) begin
		AssumePrime = 1;
	end	else if (num==16'd7253) begin
		AssumePrime = 1;
	end	else if (num==16'd7283) begin
		AssumePrime = 1;
	end	else if (num==16'd7297) begin
		AssumePrime = 1;
	end	else if (num==16'd7307) begin
		AssumePrime = 1;
	end	else if (num==16'd7309) begin
		AssumePrime = 1;
	end	else if (num==16'd7321) begin
		AssumePrime = 1;
	end	else if (num==16'd7331) begin
		AssumePrime = 1;
	end	else if (num==16'd7333) begin
		AssumePrime = 1;
	end	else if (num==16'd7349) begin
		AssumePrime = 1;
	end	else if (num==16'd7351) begin
		AssumePrime = 1;
	end	else if (num==16'd7369) begin
		AssumePrime = 1;
	end	else if (num==16'd7393) begin
		AssumePrime = 1;
	end	else if (num==16'd7411) begin
		AssumePrime = 1;
	end	else if (num==16'd7417) begin
		AssumePrime = 1;
	end	else if (num==16'd7433) begin
		AssumePrime = 1;
	end	else if (num==16'd7451) begin
		AssumePrime = 1;
	end	else if (num==16'd7457) begin
		AssumePrime = 1;
	end	else if (num==16'd7459) begin
		AssumePrime = 1;
	end	else if (num==16'd7477) begin
		AssumePrime = 1;
	end	else if (num==16'd7481) begin
		AssumePrime = 1;
	end	else if (num==16'd7487) begin
		AssumePrime = 1;
	end	else if (num==16'd7489) begin
		AssumePrime = 1;
	end	else if (num==16'd7499) begin
		AssumePrime = 1;
	end	else if (num==16'd7507) begin
		AssumePrime = 1;
	end	else if (num==16'd7517) begin
		AssumePrime = 1;
	end	else if (num==16'd7523) begin
		AssumePrime = 1;
	end	else if (num==16'd7529) begin
		AssumePrime = 1;
	end	else if (num==16'd7537) begin
		AssumePrime = 1;
	end	else if (num==16'd7541) begin
		AssumePrime = 1;
	end	else if (num==16'd7547) begin
		AssumePrime = 1;
	end	else if (num==16'd7549) begin
		AssumePrime = 1;
	end	else if (num==16'd7559) begin
		AssumePrime = 1;
	end	else if (num==16'd7561) begin
		AssumePrime = 1;
	end	else if (num==16'd7573) begin
		AssumePrime = 1;
	end	else if (num==16'd7577) begin
		AssumePrime = 1;
	end	else if (num==16'd7583) begin
		AssumePrime = 1;
	end	else if (num==16'd7589) begin
		AssumePrime = 1;
	end	else if (num==16'd7591) begin
		AssumePrime = 1;
	end	else if (num==16'd7603) begin
		AssumePrime = 1;
	end	else if (num==16'd7607) begin
		AssumePrime = 1;
	end	else if (num==16'd7621) begin
		AssumePrime = 1;
	end	else if (num==16'd7639) begin
		AssumePrime = 1;
	end	else if (num==16'd7643) begin
		AssumePrime = 1;
	end	else if (num==16'd7649) begin
		AssumePrime = 1;
	end	else if (num==16'd7669) begin
		AssumePrime = 1;
	end	else if (num==16'd7673) begin
		AssumePrime = 1;
	end	else if (num==16'd7681) begin
		AssumePrime = 1;
	end	else if (num==16'd7687) begin
		AssumePrime = 1;
	end	else if (num==16'd7691) begin
		AssumePrime = 1;
	end	else if (num==16'd7699) begin
		AssumePrime = 1;
	end	else if (num==16'd7703) begin
		AssumePrime = 1;
	end	else if (num==16'd7717) begin
		AssumePrime = 1;
	end	else if (num==16'd7723) begin
		AssumePrime = 1;
	end	else if (num==16'd7727) begin
		AssumePrime = 1;
	end	else if (num==16'd7741) begin
		AssumePrime = 1;
	end	else if (num==16'd7753) begin
		AssumePrime = 1;
	end	else if (num==16'd7757) begin
		AssumePrime = 1;
	end	else if (num==16'd7759) begin
		AssumePrime = 1;
	end	else if (num==16'd7789) begin
		AssumePrime = 1;
	end	else if (num==16'd7793) begin
		AssumePrime = 1;
	end	else if (num==16'd7817) begin
		AssumePrime = 1;
	end	else if (num==16'd7823) begin
		AssumePrime = 1;
	end	else if (num==16'd7829) begin
		AssumePrime = 1;
	end	else if (num==16'd7841) begin
		AssumePrime = 1;
	end	else if (num==16'd7853) begin
		AssumePrime = 1;
	end	else if (num==16'd7867) begin
		AssumePrime = 1;
	end	else if (num==16'd7873) begin
		AssumePrime = 1;
	end	else if (num==16'd7877) begin
		AssumePrime = 1;
	end	else if (num==16'd7879) begin
		AssumePrime = 1;
	end	else if (num==16'd7883) begin
		AssumePrime = 1;
	end	else if (num==16'd7901) begin
		AssumePrime = 1;
	end	else if (num==16'd7907) begin
		AssumePrime = 1;
	end	else if (num==16'd7919) begin
		AssumePrime = 1;
	end	else if (num==16'd7927) begin
		AssumePrime = 1;
	end	else if (num==16'd7933) begin
		AssumePrime = 1;
	end	else if (num==16'd7937) begin
		AssumePrime = 1;
	end	else if (num==16'd7949) begin
		AssumePrime = 1;
	end	else if (num==16'd7951) begin
		AssumePrime = 1;
	end	else if (num==16'd7963) begin
		AssumePrime = 1;
	end	else if (num==16'd7993) begin
		AssumePrime = 1;
	end	else if (num==16'd8009) begin
		AssumePrime = 1;
	end	else if (num==16'd8011) begin
		AssumePrime = 1;
	end	else if (num==16'd8017) begin
		AssumePrime = 1;
	end	else if (num==16'd8039) begin
		AssumePrime = 1;
	end	else if (num==16'd8053) begin
		AssumePrime = 1;
	end	else if (num==16'd8059) begin
		AssumePrime = 1;
	end	else if (num==16'd8069) begin
		AssumePrime = 1;
	end	else if (num==16'd8081) begin
		AssumePrime = 1;
	end	else if (num==16'd8087) begin
		AssumePrime = 1;
	end	else if (num==16'd8089) begin
		AssumePrime = 1;
	end	else if (num==16'd8093) begin
		AssumePrime = 1;
	end	else if (num==16'd8101) begin
		AssumePrime = 1;
	end	else if (num==16'd8111) begin
		AssumePrime = 1;
	end	else if (num==16'd8117) begin
		AssumePrime = 1;
	end	else if (num==16'd8123) begin
		AssumePrime = 1;
	end	else if (num==16'd8147) begin
		AssumePrime = 1;
	end	else if (num==16'd8161) begin
		AssumePrime = 1;
	end	else if (num==16'd8167) begin
		AssumePrime = 1;
	end	else if (num==16'd8171) begin
		AssumePrime = 1;
	end	else if (num==16'd8179) begin
		AssumePrime = 1;
	end	else if (num==16'd8191) begin
		AssumePrime = 1;
	end	else if (num==16'd8209) begin
		AssumePrime = 1;
	end	else if (num==16'd8219) begin
		AssumePrime = 1;
	end	else if (num==16'd8221) begin
		AssumePrime = 1;
	end	else if (num==16'd8231) begin
		AssumePrime = 1;
	end	else if (num==16'd8233) begin
		AssumePrime = 1;
	end	else if (num==16'd8237) begin
		AssumePrime = 1;
	end	else if (num==16'd8243) begin
		AssumePrime = 1;
	end	else if (num==16'd8263) begin
		AssumePrime = 1;
	end	else if (num==16'd8269) begin
		AssumePrime = 1;
	end	else if (num==16'd8273) begin
		AssumePrime = 1;
	end	else if (num==16'd8287) begin
		AssumePrime = 1;
	end	else if (num==16'd8291) begin
		AssumePrime = 1;
	end	else if (num==16'd8293) begin
		AssumePrime = 1;
	end	else if (num==16'd8297) begin
		AssumePrime = 1;
	end	else if (num==16'd8311) begin
		AssumePrime = 1;
	end	else if (num==16'd8317) begin
		AssumePrime = 1;
	end	else if (num==16'd8329) begin
		AssumePrime = 1;
	end	else if (num==16'd8353) begin
		AssumePrime = 1;
	end	else if (num==16'd8363) begin
		AssumePrime = 1;
	end	else if (num==16'd8369) begin
		AssumePrime = 1;
	end	else if (num==16'd8377) begin
		AssumePrime = 1;
	end	else if (num==16'd8387) begin
		AssumePrime = 1;
	end	else if (num==16'd8389) begin
		AssumePrime = 1;
	end	else if (num==16'd8419) begin
		AssumePrime = 1;
	end	else if (num==16'd8423) begin
		AssumePrime = 1;
	end	else if (num==16'd8429) begin
		AssumePrime = 1;
	end	else if (num==16'd8431) begin
		AssumePrime = 1;
	end	else if (num==16'd8443) begin
		AssumePrime = 1;
	end	else if (num==16'd8447) begin
		AssumePrime = 1;
	end	else if (num==16'd8461) begin
		AssumePrime = 1;
	end	else if (num==16'd8467) begin
		AssumePrime = 1;
	end	else if (num==16'd8501) begin
		AssumePrime = 1;
	end	else if (num==16'd8513) begin
		AssumePrime = 1;
	end	else if (num==16'd8521) begin
		AssumePrime = 1;
	end	else if (num==16'd8527) begin
		AssumePrime = 1;
	end	else if (num==16'd8537) begin
		AssumePrime = 1;
	end	else if (num==16'd8539) begin
		AssumePrime = 1;
	end	else if (num==16'd8543) begin
		AssumePrime = 1;
	end	else if (num==16'd8563) begin
		AssumePrime = 1;
	end	else if (num==16'd8573) begin
		AssumePrime = 1;
	end	else if (num==16'd8581) begin
		AssumePrime = 1;
	end	else if (num==16'd8597) begin
		AssumePrime = 1;
	end	else if (num==16'd8599) begin
		AssumePrime = 1;
	end	else if (num==16'd8609) begin
		AssumePrime = 1;
	end	else if (num==16'd8623) begin
		AssumePrime = 1;
	end	else if (num==16'd8627) begin
		AssumePrime = 1;
	end	else if (num==16'd8629) begin
		AssumePrime = 1;
	end	else if (num==16'd8641) begin
		AssumePrime = 1;
	end	else if (num==16'd8647) begin
		AssumePrime = 1;
	end	else if (num==16'd8663) begin
		AssumePrime = 1;
	end	else if (num==16'd8669) begin
		AssumePrime = 1;
	end	else if (num==16'd8677) begin
		AssumePrime = 1;
	end	else if (num==16'd8681) begin
		AssumePrime = 1;
	end	else if (num==16'd8689) begin
		AssumePrime = 1;
	end	else if (num==16'd8693) begin
		AssumePrime = 1;
	end	else if (num==16'd8699) begin
		AssumePrime = 1;
	end	else if (num==16'd8707) begin
		AssumePrime = 1;
	end	else if (num==16'd8713) begin
		AssumePrime = 1;
	end	else if (num==16'd8719) begin
		AssumePrime = 1;
	end	else if (num==16'd8731) begin
		AssumePrime = 1;
	end	else if (num==16'd8737) begin
		AssumePrime = 1;
	end	else if (num==16'd8741) begin
		AssumePrime = 1;
	end	else if (num==16'd8747) begin
		AssumePrime = 1;
	end	else if (num==16'd8753) begin
		AssumePrime = 1;
	end	else if (num==16'd8761) begin
		AssumePrime = 1;
	end	else if (num==16'd8779) begin
		AssumePrime = 1;
	end	else if (num==16'd8783) begin
		AssumePrime = 1;
	end	else if (num==16'd8803) begin
		AssumePrime = 1;
	end	else if (num==16'd8807) begin
		AssumePrime = 1;
	end	else if (num==16'd8819) begin
		AssumePrime = 1;
	end	else if (num==16'd8821) begin
		AssumePrime = 1;
	end	else if (num==16'd8831) begin
		AssumePrime = 1;
	end	else if (num==16'd8837) begin
		AssumePrime = 1;
	end	else if (num==16'd8839) begin
		AssumePrime = 1;
	end	else if (num==16'd8849) begin
		AssumePrime = 1;
	end	else if (num==16'd8861) begin
		AssumePrime = 1;
	end	else if (num==16'd8863) begin
		AssumePrime = 1;
	end	else if (num==16'd8867) begin
		AssumePrime = 1;
	end	else if (num==16'd8887) begin
		AssumePrime = 1;
	end	else if (num==16'd8893) begin
		AssumePrime = 1;
	end	else if (num==16'd8923) begin
		AssumePrime = 1;
	end	else if (num==16'd8929) begin
		AssumePrime = 1;
	end	else if (num==16'd8933) begin
		AssumePrime = 1;
	end	else if (num==16'd8941) begin
		AssumePrime = 1;
	end	else if (num==16'd8951) begin
		AssumePrime = 1;
	end	else if (num==16'd8963) begin
		AssumePrime = 1;
	end	else if (num==16'd8969) begin
		AssumePrime = 1;
	end	else if (num==16'd8971) begin
		AssumePrime = 1;
	end	else if (num==16'd8999) begin
		AssumePrime = 1;
	end	else if (num==16'd9001) begin
		AssumePrime = 1;
	end	else if (num==16'd9007) begin
		AssumePrime = 1;
	end	else if (num==16'd9011) begin
		AssumePrime = 1;
	end	else if (num==16'd9013) begin
		AssumePrime = 1;
	end	else if (num==16'd9029) begin
		AssumePrime = 1;
	end	else if (num==16'd9041) begin
		AssumePrime = 1;
	end	else if (num==16'd9043) begin
		AssumePrime = 1;
	end	else if (num==16'd9049) begin
		AssumePrime = 1;
	end	else if (num==16'd9059) begin
		AssumePrime = 1;
	end	else if (num==16'd9067) begin
		AssumePrime = 1;
	end	else if (num==16'd9091) begin
		AssumePrime = 1;
	end	else if (num==16'd9103) begin
		AssumePrime = 1;
	end	else if (num==16'd9109) begin
		AssumePrime = 1;
	end	else if (num==16'd9127) begin
		AssumePrime = 1;
	end	else if (num==16'd9133) begin
		AssumePrime = 1;
	end	else if (num==16'd9137) begin
		AssumePrime = 1;
	end	else if (num==16'd9151) begin
		AssumePrime = 1;
	end	else if (num==16'd9157) begin
		AssumePrime = 1;
	end	else if (num==16'd9161) begin
		AssumePrime = 1;
	end	else if (num==16'd9173) begin
		AssumePrime = 1;
	end	else if (num==16'd9181) begin
		AssumePrime = 1;
	end	else if (num==16'd9187) begin
		AssumePrime = 1;
	end	else if (num==16'd9199) begin
		AssumePrime = 1;
	end	else if (num==16'd9203) begin
		AssumePrime = 1;
	end	else if (num==16'd9209) begin
		AssumePrime = 1;
	end	else if (num==16'd9221) begin
		AssumePrime = 1;
	end	else if (num==16'd9227) begin
		AssumePrime = 1;
	end	else if (num==16'd9239) begin
		AssumePrime = 1;
	end	else if (num==16'd9241) begin
		AssumePrime = 1;
	end	else if (num==16'd9257) begin
		AssumePrime = 1;
	end	else if (num==16'd9277) begin
		AssumePrime = 1;
	end	else if (num==16'd9281) begin
		AssumePrime = 1;
	end	else if (num==16'd9283) begin
		AssumePrime = 1;
	end	else if (num==16'd9293) begin
		AssumePrime = 1;
	end	else if (num==16'd9311) begin
		AssumePrime = 1;
	end	else if (num==16'd9319) begin
		AssumePrime = 1;
	end	else if (num==16'd9323) begin
		AssumePrime = 1;
	end	else if (num==16'd9337) begin
		AssumePrime = 1;
	end	else if (num==16'd9341) begin
		AssumePrime = 1;
	end	else if (num==16'd9343) begin
		AssumePrime = 1;
	end	else if (num==16'd9349) begin
		AssumePrime = 1;
	end	else if (num==16'd9371) begin
		AssumePrime = 1;
	end	else if (num==16'd9377) begin
		AssumePrime = 1;
	end	else if (num==16'd9391) begin
		AssumePrime = 1;
	end	else if (num==16'd9397) begin
		AssumePrime = 1;
	end	else if (num==16'd9403) begin
		AssumePrime = 1;
	end	else if (num==16'd9413) begin
		AssumePrime = 1;
	end	else if (num==16'd9419) begin
		AssumePrime = 1;
	end	else if (num==16'd9421) begin
		AssumePrime = 1;
	end	else if (num==16'd9431) begin
		AssumePrime = 1;
	end	else if (num==16'd9433) begin
		AssumePrime = 1;
	end	else if (num==16'd9437) begin
		AssumePrime = 1;
	end	else if (num==16'd9439) begin
		AssumePrime = 1;
	end	else if (num==16'd9461) begin
		AssumePrime = 1;
	end	else if (num==16'd9463) begin
		AssumePrime = 1;
	end	else if (num==16'd9467) begin
		AssumePrime = 1;
	end	else if (num==16'd9473) begin
		AssumePrime = 1;
	end	else if (num==16'd9479) begin
		AssumePrime = 1;
	end	else if (num==16'd9491) begin
		AssumePrime = 1;
	end	else if (num==16'd9497) begin
		AssumePrime = 1;
	end	else if (num==16'd9511) begin
		AssumePrime = 1;
	end	else if (num==16'd9521) begin
		AssumePrime = 1;
	end	else if (num==16'd9533) begin
		AssumePrime = 1;
	end	else if (num==16'd9539) begin
		AssumePrime = 1;
	end	else if (num==16'd9547) begin
		AssumePrime = 1;
	end	else if (num==16'd9551) begin
		AssumePrime = 1;
	end	else if (num==16'd9587) begin
		AssumePrime = 1;
	end	else if (num==16'd9601) begin
		AssumePrime = 1;
	end	else if (num==16'd9613) begin
		AssumePrime = 1;
	end	else if (num==16'd9619) begin
		AssumePrime = 1;
	end	else if (num==16'd9623) begin
		AssumePrime = 1;
	end	else if (num==16'd9629) begin
		AssumePrime = 1;
	end	else if (num==16'd9631) begin
		AssumePrime = 1;
	end	else if (num==16'd9643) begin
		AssumePrime = 1;
	end	else if (num==16'd9649) begin
		AssumePrime = 1;
	end	else if (num==16'd9661) begin
		AssumePrime = 1;
	end	else if (num==16'd9677) begin
		AssumePrime = 1;
	end	else if (num==16'd9679) begin
		AssumePrime = 1;
	end	else if (num==16'd9689) begin
		AssumePrime = 1;
	end	else if (num==16'd9697) begin
		AssumePrime = 1;
	end	else if (num==16'd9719) begin
		AssumePrime = 1;
	end	else if (num==16'd9721) begin
		AssumePrime = 1;
	end	else if (num==16'd9733) begin
		AssumePrime = 1;
	end	else if (num==16'd9739) begin
		AssumePrime = 1;
	end	else if (num==16'd9743) begin
		AssumePrime = 1;
	end	else if (num==16'd9749) begin
		AssumePrime = 1;
	end	else if (num==16'd9767) begin
		AssumePrime = 1;
	end	else if (num==16'd9769) begin
		AssumePrime = 1;
	end	else if (num==16'd9781) begin
		AssumePrime = 1;
	end	else if (num==16'd9787) begin
		AssumePrime = 1;
	end	else if (num==16'd9791) begin
		AssumePrime = 1;
	end	else if (num==16'd9803) begin
		AssumePrime = 1;
	end	else if (num==16'd9811) begin
		AssumePrime = 1;
	end	else if (num==16'd9817) begin
		AssumePrime = 1;
	end	else if (num==16'd9829) begin
		AssumePrime = 1;
	end	else if (num==16'd9833) begin
		AssumePrime = 1;
	end	else if (num==16'd9839) begin
		AssumePrime = 1;
	end	else if (num==16'd9851) begin
		AssumePrime = 1;
	end	else if (num==16'd9857) begin
		AssumePrime = 1;
	end	else if (num==16'd9859) begin
		AssumePrime = 1;
	end	else if (num==16'd9871) begin
		AssumePrime = 1;
	end	else if (num==16'd9883) begin
		AssumePrime = 1;
	end	else if (num==16'd9887) begin
		AssumePrime = 1;
	end	else if (num==16'd9901) begin
		AssumePrime = 1;
	end	else if (num==16'd9907) begin
		AssumePrime = 1;
	end	else if (num==16'd9923) begin
		AssumePrime = 1;
	end	else if (num==16'd9929) begin
		AssumePrime = 1;
	end	else if (num==16'd9931) begin
		AssumePrime = 1;
	end	else if (num==16'd9941) begin
		AssumePrime = 1;
	end	else if (num==16'd9949) begin
		AssumePrime = 1;
	end	else if (num==16'd9967) begin
		AssumePrime = 1;
	end	else if (num==16'd9973) begin
		AssumePrime = 1;
	end	else if (num==16'd10007) begin
		AssumePrime = 1;
	end	else if (num==16'd10009) begin
		AssumePrime = 1;
	end	else if (num==16'd10037) begin
		AssumePrime = 1;
	end	else if (num==16'd10039) begin
		AssumePrime = 1;
	end	else if (num==16'd10061) begin
		AssumePrime = 1;
	end	else if (num==16'd10067) begin
		AssumePrime = 1;
	end	else if (num==16'd10069) begin
		AssumePrime = 1;
	end	else if (num==16'd10079) begin
		AssumePrime = 1;
	end	else if (num==16'd10091) begin
		AssumePrime = 1;
	end	else if (num==16'd10093) begin
		AssumePrime = 1;
	end	else if (num==16'd10099) begin
		AssumePrime = 1;
	end	else if (num==16'd10103) begin
		AssumePrime = 1;
	end	else if (num==16'd10111) begin
		AssumePrime = 1;
	end	else if (num==16'd10133) begin
		AssumePrime = 1;
	end	else if (num==16'd10139) begin
		AssumePrime = 1;
	end	else if (num==16'd10141) begin
		AssumePrime = 1;
	end	else if (num==16'd10151) begin
		AssumePrime = 1;
	end	else if (num==16'd10159) begin
		AssumePrime = 1;
	end	else if (num==16'd10163) begin
		AssumePrime = 1;
	end	else if (num==16'd10169) begin
		AssumePrime = 1;
	end	else if (num==16'd10177) begin
		AssumePrime = 1;
	end	else if (num==16'd10181) begin
		AssumePrime = 1;
	end	else if (num==16'd10193) begin
		AssumePrime = 1;
	end	else if (num==16'd10211) begin
		AssumePrime = 1;
	end	else if (num==16'd10223) begin
		AssumePrime = 1;
	end	else if (num==16'd10243) begin
		AssumePrime = 1;
	end	else if (num==16'd10247) begin
		AssumePrime = 1;
	end	else if (num==16'd10253) begin
		AssumePrime = 1;
	end	else if (num==16'd10259) begin
		AssumePrime = 1;
	end	else if (num==16'd10267) begin
		AssumePrime = 1;
	end	else if (num==16'd10271) begin
		AssumePrime = 1;
	end	else if (num==16'd10273) begin
		AssumePrime = 1;
	end	else if (num==16'd10289) begin
		AssumePrime = 1;
	end	else if (num==16'd10301) begin
		AssumePrime = 1;
	end	else if (num==16'd10303) begin
		AssumePrime = 1;
	end	else if (num==16'd10313) begin
		AssumePrime = 1;
	end	else if (num==16'd10321) begin
		AssumePrime = 1;
	end	else if (num==16'd10331) begin
		AssumePrime = 1;
	end	else if (num==16'd10333) begin
		AssumePrime = 1;
	end	else if (num==16'd10337) begin
		AssumePrime = 1;
	end	else if (num==16'd10343) begin
		AssumePrime = 1;
	end	else if (num==16'd10357) begin
		AssumePrime = 1;
	end	else if (num==16'd10369) begin
		AssumePrime = 1;
	end	else if (num==16'd10391) begin
		AssumePrime = 1;
	end	else if (num==16'd10399) begin
		AssumePrime = 1;
	end	else if (num==16'd10427) begin
		AssumePrime = 1;
	end	else if (num==16'd10429) begin
		AssumePrime = 1;
	end	else if (num==16'd10433) begin
		AssumePrime = 1;
	end	else if (num==16'd10453) begin
		AssumePrime = 1;
	end	else if (num==16'd10457) begin
		AssumePrime = 1;
	end	else if (num==16'd10459) begin
		AssumePrime = 1;
	end	else if (num==16'd10463) begin
		AssumePrime = 1;
	end	else if (num==16'd10477) begin
		AssumePrime = 1;
	end	else if (num==16'd10487) begin
		AssumePrime = 1;
	end	else if (num==16'd10499) begin
		AssumePrime = 1;
	end	else if (num==16'd10501) begin
		AssumePrime = 1;
	end	else if (num==16'd10513) begin
		AssumePrime = 1;
	end	else if (num==16'd10529) begin
		AssumePrime = 1;
	end	else if (num==16'd10531) begin
		AssumePrime = 1;
	end	else if (num==16'd10559) begin
		AssumePrime = 1;
	end	else if (num==16'd10567) begin
		AssumePrime = 1;
	end	else if (num==16'd10589) begin
		AssumePrime = 1;
	end	else if (num==16'd10597) begin
		AssumePrime = 1;
	end	else if (num==16'd10601) begin
		AssumePrime = 1;
	end	else if (num==16'd10607) begin
		AssumePrime = 1;
	end	else if (num==16'd10613) begin
		AssumePrime = 1;
	end	else if (num==16'd10627) begin
		AssumePrime = 1;
	end	else if (num==16'd10631) begin
		AssumePrime = 1;
	end	else if (num==16'd10639) begin
		AssumePrime = 1;
	end	else if (num==16'd10651) begin
		AssumePrime = 1;
	end	else if (num==16'd10657) begin
		AssumePrime = 1;
	end	else if (num==16'd10663) begin
		AssumePrime = 1;
	end	else if (num==16'd10667) begin
		AssumePrime = 1;
	end	else if (num==16'd10687) begin
		AssumePrime = 1;
	end	else if (num==16'd10691) begin
		AssumePrime = 1;
	end	else if (num==16'd10709) begin
		AssumePrime = 1;
	end	else if (num==16'd10711) begin
		AssumePrime = 1;
	end	else if (num==16'd10723) begin
		AssumePrime = 1;
	end	else if (num==16'd10729) begin
		AssumePrime = 1;
	end	else if (num==16'd10733) begin
		AssumePrime = 1;
	end	else if (num==16'd10739) begin
		AssumePrime = 1;
	end	else if (num==16'd10753) begin
		AssumePrime = 1;
	end	else if (num==16'd10771) begin
		AssumePrime = 1;
	end	else if (num==16'd10781) begin
		AssumePrime = 1;
	end	else if (num==16'd10789) begin
		AssumePrime = 1;
	end	else if (num==16'd10799) begin
		AssumePrime = 1;
	end	else if (num==16'd10831) begin
		AssumePrime = 1;
	end	else if (num==16'd10837) begin
		AssumePrime = 1;
	end	else if (num==16'd10847) begin
		AssumePrime = 1;
	end	else if (num==16'd10853) begin
		AssumePrime = 1;
	end	else if (num==16'd10859) begin
		AssumePrime = 1;
	end	else if (num==16'd10861) begin
		AssumePrime = 1;
	end	else if (num==16'd10867) begin
		AssumePrime = 1;
	end	else if (num==16'd10883) begin
		AssumePrime = 1;
	end	else if (num==16'd10889) begin
		AssumePrime = 1;
	end	else if (num==16'd10891) begin
		AssumePrime = 1;
	end	else if (num==16'd10903) begin
		AssumePrime = 1;
	end	else if (num==16'd10909) begin
		AssumePrime = 1;
	end	else if (num==16'd10937) begin
		AssumePrime = 1;
	end	else if (num==16'd10939) begin
		AssumePrime = 1;
	end	else if (num==16'd10949) begin
		AssumePrime = 1;
	end	else if (num==16'd10957) begin
		AssumePrime = 1;
	end	else if (num==16'd10973) begin
		AssumePrime = 1;
	end	else if (num==16'd10979) begin
		AssumePrime = 1;
	end	else if (num==16'd10987) begin
		AssumePrime = 1;
	end	else if (num==16'd10993) begin
		AssumePrime = 1;
	end	else if (num==16'd11003) begin
		AssumePrime = 1;
	end	else if (num==16'd11027) begin
		AssumePrime = 1;
	end	else if (num==16'd11047) begin
		AssumePrime = 1;
	end	else if (num==16'd11057) begin
		AssumePrime = 1;
	end	else if (num==16'd11059) begin
		AssumePrime = 1;
	end	else if (num==16'd11069) begin
		AssumePrime = 1;
	end	else if (num==16'd11071) begin
		AssumePrime = 1;
	end	else if (num==16'd11083) begin
		AssumePrime = 1;
	end	else if (num==16'd11087) begin
		AssumePrime = 1;
	end	else if (num==16'd11093) begin
		AssumePrime = 1;
	end	else if (num==16'd11113) begin
		AssumePrime = 1;
	end	else if (num==16'd11117) begin
		AssumePrime = 1;
	end	else if (num==16'd11119) begin
		AssumePrime = 1;
	end	else if (num==16'd11131) begin
		AssumePrime = 1;
	end	else if (num==16'd11149) begin
		AssumePrime = 1;
	end	else if (num==16'd11159) begin
		AssumePrime = 1;
	end	else if (num==16'd11161) begin
		AssumePrime = 1;
	end	else if (num==16'd11171) begin
		AssumePrime = 1;
	end	else if (num==16'd11173) begin
		AssumePrime = 1;
	end	else if (num==16'd11177) begin
		AssumePrime = 1;
	end	else if (num==16'd11197) begin
		AssumePrime = 1;
	end	else if (num==16'd11213) begin
		AssumePrime = 1;
	end	else if (num==16'd11239) begin
		AssumePrime = 1;
	end	else if (num==16'd11243) begin
		AssumePrime = 1;
	end	else if (num==16'd11251) begin
		AssumePrime = 1;
	end	else if (num==16'd11257) begin
		AssumePrime = 1;
	end	else if (num==16'd11261) begin
		AssumePrime = 1;
	end	else if (num==16'd11273) begin
		AssumePrime = 1;
	end	else if (num==16'd11279) begin
		AssumePrime = 1;
	end	else if (num==16'd11287) begin
		AssumePrime = 1;
	end	else if (num==16'd11299) begin
		AssumePrime = 1;
	end	else if (num==16'd11311) begin
		AssumePrime = 1;
	end	else if (num==16'd11317) begin
		AssumePrime = 1;
	end	else if (num==16'd11321) begin
		AssumePrime = 1;
	end	else if (num==16'd11329) begin
		AssumePrime = 1;
	end	else if (num==16'd11351) begin
		AssumePrime = 1;
	end	else if (num==16'd11353) begin
		AssumePrime = 1;
	end	else if (num==16'd11369) begin
		AssumePrime = 1;
	end	else if (num==16'd11383) begin
		AssumePrime = 1;
	end	else if (num==16'd11393) begin
		AssumePrime = 1;
	end	else if (num==16'd11399) begin
		AssumePrime = 1;
	end	else if (num==16'd11411) begin
		AssumePrime = 1;
	end	else if (num==16'd11423) begin
		AssumePrime = 1;
	end	else if (num==16'd11437) begin
		AssumePrime = 1;
	end	else if (num==16'd11443) begin
		AssumePrime = 1;
	end	else if (num==16'd11447) begin
		AssumePrime = 1;
	end	else if (num==16'd11467) begin
		AssumePrime = 1;
	end	else if (num==16'd11471) begin
		AssumePrime = 1;
	end	else if (num==16'd11483) begin
		AssumePrime = 1;
	end	else if (num==16'd11489) begin
		AssumePrime = 1;
	end	else if (num==16'd11491) begin
		AssumePrime = 1;
	end	else if (num==16'd11497) begin
		AssumePrime = 1;
	end	else if (num==16'd11503) begin
		AssumePrime = 1;
	end	else if (num==16'd11519) begin
		AssumePrime = 1;
	end	else if (num==16'd11527) begin
		AssumePrime = 1;
	end	else if (num==16'd11549) begin
		AssumePrime = 1;
	end	else if (num==16'd11551) begin
		AssumePrime = 1;
	end	else if (num==16'd11579) begin
		AssumePrime = 1;
	end	else if (num==16'd11587) begin
		AssumePrime = 1;
	end	else if (num==16'd11593) begin
		AssumePrime = 1;
	end	else if (num==16'd11597) begin
		AssumePrime = 1;
	end	else if (num==16'd11617) begin
		AssumePrime = 1;
	end	else if (num==16'd11621) begin
		AssumePrime = 1;
	end	else if (num==16'd11633) begin
		AssumePrime = 1;
	end	else if (num==16'd11657) begin
		AssumePrime = 1;
	end	else if (num==16'd11677) begin
		AssumePrime = 1;
	end	else if (num==16'd11681) begin
		AssumePrime = 1;
	end	else if (num==16'd11689) begin
		AssumePrime = 1;
	end	else if (num==16'd11699) begin
		AssumePrime = 1;
	end	else if (num==16'd11701) begin
		AssumePrime = 1;
	end	else if (num==16'd11717) begin
		AssumePrime = 1;
	end	else if (num==16'd11719) begin
		AssumePrime = 1;
	end	else if (num==16'd11731) begin
		AssumePrime = 1;
	end	else if (num==16'd11743) begin
		AssumePrime = 1;
	end	else if (num==16'd11777) begin
		AssumePrime = 1;
	end	else if (num==16'd11779) begin
		AssumePrime = 1;
	end	else if (num==16'd11783) begin
		AssumePrime = 1;
	end	else if (num==16'd11789) begin
		AssumePrime = 1;
	end	else if (num==16'd11801) begin
		AssumePrime = 1;
	end	else if (num==16'd11807) begin
		AssumePrime = 1;
	end	else if (num==16'd11813) begin
		AssumePrime = 1;
	end	else if (num==16'd11821) begin
		AssumePrime = 1;
	end	else if (num==16'd11827) begin
		AssumePrime = 1;
	end	else if (num==16'd11831) begin
		AssumePrime = 1;
	end	else if (num==16'd11833) begin
		AssumePrime = 1;
	end	else if (num==16'd11839) begin
		AssumePrime = 1;
	end	else if (num==16'd11863) begin
		AssumePrime = 1;
	end	else if (num==16'd11867) begin
		AssumePrime = 1;
	end	else if (num==16'd11887) begin
		AssumePrime = 1;
	end	else if (num==16'd11897) begin
		AssumePrime = 1;
	end	else if (num==16'd11903) begin
		AssumePrime = 1;
	end	else if (num==16'd11909) begin
		AssumePrime = 1;
	end	else if (num==16'd11923) begin
		AssumePrime = 1;
	end	else if (num==16'd11927) begin
		AssumePrime = 1;
	end	else if (num==16'd11933) begin
		AssumePrime = 1;
	end	else if (num==16'd11939) begin
		AssumePrime = 1;
	end	else if (num==16'd11941) begin
		AssumePrime = 1;
	end	else if (num==16'd11953) begin
		AssumePrime = 1;
	end	else if (num==16'd11959) begin
		AssumePrime = 1;
	end	else if (num==16'd11969) begin
		AssumePrime = 1;
	end	else if (num==16'd11971) begin
		AssumePrime = 1;
	end	else if (num==16'd11981) begin
		AssumePrime = 1;
	end	else if (num==16'd11987) begin
		AssumePrime = 1;
	end	else if (num==16'd12007) begin
		AssumePrime = 1;
	end	else if (num==16'd12011) begin
		AssumePrime = 1;
	end	else if (num==16'd12037) begin
		AssumePrime = 1;
	end	else if (num==16'd12041) begin
		AssumePrime = 1;
	end	else if (num==16'd12043) begin
		AssumePrime = 1;
	end	else if (num==16'd12049) begin
		AssumePrime = 1;
	end	else if (num==16'd12071) begin
		AssumePrime = 1;
	end	else if (num==16'd12073) begin
		AssumePrime = 1;
	end	else if (num==16'd12097) begin
		AssumePrime = 1;
	end	else if (num==16'd12101) begin
		AssumePrime = 1;
	end	else if (num==16'd12107) begin
		AssumePrime = 1;
	end	else if (num==16'd12109) begin
		AssumePrime = 1;
	end	else if (num==16'd12113) begin
		AssumePrime = 1;
	end	else if (num==16'd12119) begin
		AssumePrime = 1;
	end	else if (num==16'd12143) begin
		AssumePrime = 1;
	end	else if (num==16'd12149) begin
		AssumePrime = 1;
	end	else if (num==16'd12157) begin
		AssumePrime = 1;
	end	else if (num==16'd12161) begin
		AssumePrime = 1;
	end	else if (num==16'd12163) begin
		AssumePrime = 1;
	end	else if (num==16'd12197) begin
		AssumePrime = 1;
	end	else if (num==16'd12203) begin
		AssumePrime = 1;
	end	else if (num==16'd12211) begin
		AssumePrime = 1;
	end	else if (num==16'd12227) begin
		AssumePrime = 1;
	end	else if (num==16'd12239) begin
		AssumePrime = 1;
	end	else if (num==16'd12241) begin
		AssumePrime = 1;
	end	else if (num==16'd12251) begin
		AssumePrime = 1;
	end	else if (num==16'd12253) begin
		AssumePrime = 1;
	end	else if (num==16'd12263) begin
		AssumePrime = 1;
	end	else if (num==16'd12269) begin
		AssumePrime = 1;
	end	else if (num==16'd12277) begin
		AssumePrime = 1;
	end	else if (num==16'd12281) begin
		AssumePrime = 1;
	end	else if (num==16'd12289) begin
		AssumePrime = 1;
	end	else if (num==16'd12301) begin
		AssumePrime = 1;
	end	else if (num==16'd12323) begin
		AssumePrime = 1;
	end	else if (num==16'd12329) begin
		AssumePrime = 1;
	end	else if (num==16'd12343) begin
		AssumePrime = 1;
	end	else if (num==16'd12347) begin
		AssumePrime = 1;
	end	else if (num==16'd12373) begin
		AssumePrime = 1;
	end	else if (num==16'd12377) begin
		AssumePrime = 1;
	end	else if (num==16'd12379) begin
		AssumePrime = 1;
	end	else if (num==16'd12391) begin
		AssumePrime = 1;
	end	else if (num==16'd12401) begin
		AssumePrime = 1;
	end	else if (num==16'd12409) begin
		AssumePrime = 1;
	end	else if (num==16'd12413) begin
		AssumePrime = 1;
	end	else if (num==16'd12421) begin
		AssumePrime = 1;
	end	else if (num==16'd12433) begin
		AssumePrime = 1;
	end	else if (num==16'd12437) begin
		AssumePrime = 1;
	end	else if (num==16'd12451) begin
		AssumePrime = 1;
	end	else if (num==16'd12457) begin
		AssumePrime = 1;
	end	else if (num==16'd12473) begin
		AssumePrime = 1;
	end	else if (num==16'd12479) begin
		AssumePrime = 1;
	end	else if (num==16'd12487) begin
		AssumePrime = 1;
	end	else if (num==16'd12491) begin
		AssumePrime = 1;
	end	else if (num==16'd12497) begin
		AssumePrime = 1;
	end	else if (num==16'd12503) begin
		AssumePrime = 1;
	end	else if (num==16'd12511) begin
		AssumePrime = 1;
	end	else if (num==16'd12517) begin
		AssumePrime = 1;
	end	else if (num==16'd12527) begin
		AssumePrime = 1;
	end	else if (num==16'd12539) begin
		AssumePrime = 1;
	end	else if (num==16'd12541) begin
		AssumePrime = 1;
	end	else if (num==16'd12547) begin
		AssumePrime = 1;
	end	else if (num==16'd12553) begin
		AssumePrime = 1;
	end	else if (num==16'd12569) begin
		AssumePrime = 1;
	end	else if (num==16'd12577) begin
		AssumePrime = 1;
	end	else if (num==16'd12583) begin
		AssumePrime = 1;
	end	else if (num==16'd12589) begin
		AssumePrime = 1;
	end	else if (num==16'd12601) begin
		AssumePrime = 1;
	end	else if (num==16'd12611) begin
		AssumePrime = 1;
	end	else if (num==16'd12613) begin
		AssumePrime = 1;
	end	else if (num==16'd12619) begin
		AssumePrime = 1;
	end	else if (num==16'd12637) begin
		AssumePrime = 1;
	end	else if (num==16'd12641) begin
		AssumePrime = 1;
	end	else if (num==16'd12647) begin
		AssumePrime = 1;
	end	else if (num==16'd12653) begin
		AssumePrime = 1;
	end	else if (num==16'd12659) begin
		AssumePrime = 1;
	end	else if (num==16'd12671) begin
		AssumePrime = 1;
	end	else if (num==16'd12689) begin
		AssumePrime = 1;
	end	else if (num==16'd12697) begin
		AssumePrime = 1;
	end	else if (num==16'd12703) begin
		AssumePrime = 1;
	end	else if (num==16'd12713) begin
		AssumePrime = 1;
	end	else if (num==16'd12721) begin
		AssumePrime = 1;
	end	else if (num==16'd12739) begin
		AssumePrime = 1;
	end	else if (num==16'd12743) begin
		AssumePrime = 1;
	end	else if (num==16'd12757) begin
		AssumePrime = 1;
	end	else if (num==16'd12763) begin
		AssumePrime = 1;
	end	else if (num==16'd12781) begin
		AssumePrime = 1;
	end	else if (num==16'd12791) begin
		AssumePrime = 1;
	end	else if (num==16'd12799) begin
		AssumePrime = 1;
	end	else if (num==16'd12809) begin
		AssumePrime = 1;
	end	else if (num==16'd12821) begin
		AssumePrime = 1;
	end	else if (num==16'd12823) begin
		AssumePrime = 1;
	end	else if (num==16'd12829) begin
		AssumePrime = 1;
	end	else if (num==16'd12841) begin
		AssumePrime = 1;
	end	else if (num==16'd12853) begin
		AssumePrime = 1;
	end	else if (num==16'd12889) begin
		AssumePrime = 1;
	end	else if (num==16'd12893) begin
		AssumePrime = 1;
	end	else if (num==16'd12899) begin
		AssumePrime = 1;
	end	else if (num==16'd12907) begin
		AssumePrime = 1;
	end	else if (num==16'd12911) begin
		AssumePrime = 1;
	end	else if (num==16'd12917) begin
		AssumePrime = 1;
	end	else if (num==16'd12919) begin
		AssumePrime = 1;
	end	else if (num==16'd12923) begin
		AssumePrime = 1;
	end	else if (num==16'd12941) begin
		AssumePrime = 1;
	end	else if (num==16'd12953) begin
		AssumePrime = 1;
	end	else if (num==16'd12959) begin
		AssumePrime = 1;
	end	else if (num==16'd12967) begin
		AssumePrime = 1;
	end	else if (num==16'd12973) begin
		AssumePrime = 1;
	end	else if (num==16'd12979) begin
		AssumePrime = 1;
	end	else if (num==16'd12983) begin
		AssumePrime = 1;
	end	else if (num==16'd13001) begin
		AssumePrime = 1;
	end	else if (num==16'd13003) begin
		AssumePrime = 1;
	end	else if (num==16'd13007) begin
		AssumePrime = 1;
	end	else if (num==16'd13009) begin
		AssumePrime = 1;
	end	else if (num==16'd13033) begin
		AssumePrime = 1;
	end	else if (num==16'd13037) begin
		AssumePrime = 1;
	end	else if (num==16'd13043) begin
		AssumePrime = 1;
	end	else if (num==16'd13049) begin
		AssumePrime = 1;
	end	else if (num==16'd13063) begin
		AssumePrime = 1;
	end	else if (num==16'd13093) begin
		AssumePrime = 1;
	end	else if (num==16'd13099) begin
		AssumePrime = 1;
	end	else if (num==16'd13103) begin
		AssumePrime = 1;
	end	else if (num==16'd13109) begin
		AssumePrime = 1;
	end	else if (num==16'd13121) begin
		AssumePrime = 1;
	end	else if (num==16'd13127) begin
		AssumePrime = 1;
	end	else if (num==16'd13147) begin
		AssumePrime = 1;
	end	else if (num==16'd13151) begin
		AssumePrime = 1;
	end	else if (num==16'd13159) begin
		AssumePrime = 1;
	end	else if (num==16'd13163) begin
		AssumePrime = 1;
	end	else if (num==16'd13171) begin
		AssumePrime = 1;
	end	else if (num==16'd13177) begin
		AssumePrime = 1;
	end	else if (num==16'd13183) begin
		AssumePrime = 1;
	end	else if (num==16'd13187) begin
		AssumePrime = 1;
	end	else if (num==16'd13217) begin
		AssumePrime = 1;
	end	else if (num==16'd13219) begin
		AssumePrime = 1;
	end	else if (num==16'd13229) begin
		AssumePrime = 1;
	end	else if (num==16'd13241) begin
		AssumePrime = 1;
	end	else if (num==16'd13249) begin
		AssumePrime = 1;
	end	else if (num==16'd13259) begin
		AssumePrime = 1;
	end	else if (num==16'd13267) begin
		AssumePrime = 1;
	end	else if (num==16'd13291) begin
		AssumePrime = 1;
	end	else if (num==16'd13297) begin
		AssumePrime = 1;
	end	else if (num==16'd13309) begin
		AssumePrime = 1;
	end	else if (num==16'd13313) begin
		AssumePrime = 1;
	end	else if (num==16'd13327) begin
		AssumePrime = 1;
	end	else if (num==16'd13331) begin
		AssumePrime = 1;
	end	else if (num==16'd13337) begin
		AssumePrime = 1;
	end	else if (num==16'd13339) begin
		AssumePrime = 1;
	end	else if (num==16'd13367) begin
		AssumePrime = 1;
	end	else if (num==16'd13381) begin
		AssumePrime = 1;
	end	else if (num==16'd13397) begin
		AssumePrime = 1;
	end	else if (num==16'd13399) begin
		AssumePrime = 1;
	end	else if (num==16'd13411) begin
		AssumePrime = 1;
	end	else if (num==16'd13417) begin
		AssumePrime = 1;
	end	else if (num==16'd13421) begin
		AssumePrime = 1;
	end	else if (num==16'd13441) begin
		AssumePrime = 1;
	end	else if (num==16'd13451) begin
		AssumePrime = 1;
	end	else if (num==16'd13457) begin
		AssumePrime = 1;
	end	else if (num==16'd13463) begin
		AssumePrime = 1;
	end	else if (num==16'd13469) begin
		AssumePrime = 1;
	end	else if (num==16'd13477) begin
		AssumePrime = 1;
	end	else if (num==16'd13487) begin
		AssumePrime = 1;
	end	else if (num==16'd13499) begin
		AssumePrime = 1;
	end	else if (num==16'd13513) begin
		AssumePrime = 1;
	end	else if (num==16'd13523) begin
		AssumePrime = 1;
	end	else if (num==16'd13537) begin
		AssumePrime = 1;
	end	else if (num==16'd13553) begin
		AssumePrime = 1;
	end	else if (num==16'd13567) begin
		AssumePrime = 1;
	end	else if (num==16'd13577) begin
		AssumePrime = 1;
	end	else if (num==16'd13591) begin
		AssumePrime = 1;
	end	else if (num==16'd13597) begin
		AssumePrime = 1;
	end	else if (num==16'd13613) begin
		AssumePrime = 1;
	end	else if (num==16'd13619) begin
		AssumePrime = 1;
	end	else if (num==16'd13627) begin
		AssumePrime = 1;
	end	else if (num==16'd13633) begin
		AssumePrime = 1;
	end	else if (num==16'd13649) begin
		AssumePrime = 1;
	end	else if (num==16'd13669) begin
		AssumePrime = 1;
	end	else if (num==16'd13679) begin
		AssumePrime = 1;
	end	else if (num==16'd13681) begin
		AssumePrime = 1;
	end	else if (num==16'd13687) begin
		AssumePrime = 1;
	end	else if (num==16'd13691) begin
		AssumePrime = 1;
	end	else if (num==16'd13693) begin
		AssumePrime = 1;
	end	else if (num==16'd13697) begin
		AssumePrime = 1;
	end	else if (num==16'd13709) begin
		AssumePrime = 1;
	end	else if (num==16'd13711) begin
		AssumePrime = 1;
	end	else if (num==16'd13721) begin
		AssumePrime = 1;
	end	else if (num==16'd13723) begin
		AssumePrime = 1;
	end	else if (num==16'd13729) begin
		AssumePrime = 1;
	end	else if (num==16'd13751) begin
		AssumePrime = 1;
	end	else if (num==16'd13757) begin
		AssumePrime = 1;
	end	else if (num==16'd13759) begin
		AssumePrime = 1;
	end	else if (num==16'd13763) begin
		AssumePrime = 1;
	end	else if (num==16'd13781) begin
		AssumePrime = 1;
	end	else if (num==16'd13789) begin
		AssumePrime = 1;
	end	else if (num==16'd13799) begin
		AssumePrime = 1;
	end	else if (num==16'd13807) begin
		AssumePrime = 1;
	end	else if (num==16'd13829) begin
		AssumePrime = 1;
	end	else if (num==16'd13831) begin
		AssumePrime = 1;
	end	else if (num==16'd13841) begin
		AssumePrime = 1;
	end	else if (num==16'd13859) begin
		AssumePrime = 1;
	end	else if (num==16'd13873) begin
		AssumePrime = 1;
	end	else if (num==16'd13877) begin
		AssumePrime = 1;
	end	else if (num==16'd13879) begin
		AssumePrime = 1;
	end	else if (num==16'd13883) begin
		AssumePrime = 1;
	end	else if (num==16'd13901) begin
		AssumePrime = 1;
	end	else if (num==16'd13903) begin
		AssumePrime = 1;
	end	else if (num==16'd13907) begin
		AssumePrime = 1;
	end	else if (num==16'd13913) begin
		AssumePrime = 1;
	end	else if (num==16'd13921) begin
		AssumePrime = 1;
	end	else if (num==16'd13931) begin
		AssumePrime = 1;
	end	else if (num==16'd13933) begin
		AssumePrime = 1;
	end	else if (num==16'd13963) begin
		AssumePrime = 1;
	end	else if (num==16'd13967) begin
		AssumePrime = 1;
	end	else if (num==16'd13997) begin
		AssumePrime = 1;
	end	else if (num==16'd13999) begin
		AssumePrime = 1;
	end	else if (num==16'd14009) begin
		AssumePrime = 1;
	end	else if (num==16'd14011) begin
		AssumePrime = 1;
	end	else if (num==16'd14029) begin
		AssumePrime = 1;
	end	else if (num==16'd14033) begin
		AssumePrime = 1;
	end	else if (num==16'd14051) begin
		AssumePrime = 1;
	end	else if (num==16'd14057) begin
		AssumePrime = 1;
	end	else if (num==16'd14071) begin
		AssumePrime = 1;
	end	else if (num==16'd14081) begin
		AssumePrime = 1;
	end	else if (num==16'd14083) begin
		AssumePrime = 1;
	end	else if (num==16'd14087) begin
		AssumePrime = 1;
	end	else if (num==16'd14107) begin
		AssumePrime = 1;
	end	else if (num==16'd14143) begin
		AssumePrime = 1;
	end	else if (num==16'd14149) begin
		AssumePrime = 1;
	end	else if (num==16'd14153) begin
		AssumePrime = 1;
	end	else if (num==16'd14159) begin
		AssumePrime = 1;
	end	else if (num==16'd14173) begin
		AssumePrime = 1;
	end	else if (num==16'd14177) begin
		AssumePrime = 1;
	end	else if (num==16'd14197) begin
		AssumePrime = 1;
	end	else if (num==16'd14207) begin
		AssumePrime = 1;
	end	else if (num==16'd14221) begin
		AssumePrime = 1;
	end	else if (num==16'd14243) begin
		AssumePrime = 1;
	end	else if (num==16'd14249) begin
		AssumePrime = 1;
	end	else if (num==16'd14251) begin
		AssumePrime = 1;
	end	else if (num==16'd14281) begin
		AssumePrime = 1;
	end	else if (num==16'd14293) begin
		AssumePrime = 1;
	end	else if (num==16'd14303) begin
		AssumePrime = 1;
	end	else if (num==16'd14321) begin
		AssumePrime = 1;
	end	else if (num==16'd14323) begin
		AssumePrime = 1;
	end	else if (num==16'd14327) begin
		AssumePrime = 1;
	end	else if (num==16'd14341) begin
		AssumePrime = 1;
	end	else if (num==16'd14347) begin
		AssumePrime = 1;
	end	else if (num==16'd14369) begin
		AssumePrime = 1;
	end	else if (num==16'd14387) begin
		AssumePrime = 1;
	end	else if (num==16'd14389) begin
		AssumePrime = 1;
	end	else if (num==16'd14401) begin
		AssumePrime = 1;
	end	else if (num==16'd14407) begin
		AssumePrime = 1;
	end	else if (num==16'd14411) begin
		AssumePrime = 1;
	end	else if (num==16'd14419) begin
		AssumePrime = 1;
	end	else if (num==16'd14423) begin
		AssumePrime = 1;
	end	else if (num==16'd14431) begin
		AssumePrime = 1;
	end	else if (num==16'd14437) begin
		AssumePrime = 1;
	end	else if (num==16'd14447) begin
		AssumePrime = 1;
	end	else if (num==16'd14449) begin
		AssumePrime = 1;
	end	else if (num==16'd14461) begin
		AssumePrime = 1;
	end	else if (num==16'd14479) begin
		AssumePrime = 1;
	end	else if (num==16'd14489) begin
		AssumePrime = 1;
	end	else if (num==16'd14503) begin
		AssumePrime = 1;
	end	else if (num==16'd14519) begin
		AssumePrime = 1;
	end	else if (num==16'd14533) begin
		AssumePrime = 1;
	end	else if (num==16'd14537) begin
		AssumePrime = 1;
	end	else if (num==16'd14543) begin
		AssumePrime = 1;
	end	else if (num==16'd14549) begin
		AssumePrime = 1;
	end	else if (num==16'd14551) begin
		AssumePrime = 1;
	end	else if (num==16'd14557) begin
		AssumePrime = 1;
	end	else if (num==16'd14561) begin
		AssumePrime = 1;
	end	else if (num==16'd14563) begin
		AssumePrime = 1;
	end	else if (num==16'd14591) begin
		AssumePrime = 1;
	end	else if (num==16'd14593) begin
		AssumePrime = 1;
	end	else if (num==16'd14621) begin
		AssumePrime = 1;
	end	else if (num==16'd14627) begin
		AssumePrime = 1;
	end	else if (num==16'd14629) begin
		AssumePrime = 1;
	end	else if (num==16'd14633) begin
		AssumePrime = 1;
	end	else if (num==16'd14639) begin
		AssumePrime = 1;
	end	else if (num==16'd14653) begin
		AssumePrime = 1;
	end	else if (num==16'd14657) begin
		AssumePrime = 1;
	end	else if (num==16'd14669) begin
		AssumePrime = 1;
	end	else if (num==16'd14683) begin
		AssumePrime = 1;
	end	else if (num==16'd14699) begin
		AssumePrime = 1;
	end	else if (num==16'd14713) begin
		AssumePrime = 1;
	end	else if (num==16'd14717) begin
		AssumePrime = 1;
	end	else if (num==16'd14723) begin
		AssumePrime = 1;
	end	else if (num==16'd14731) begin
		AssumePrime = 1;
	end	else if (num==16'd14737) begin
		AssumePrime = 1;
	end	else if (num==16'd14741) begin
		AssumePrime = 1;
	end	else if (num==16'd14747) begin
		AssumePrime = 1;
	end	else if (num==16'd14753) begin
		AssumePrime = 1;
	end	else if (num==16'd14759) begin
		AssumePrime = 1;
	end	else if (num==16'd14767) begin
		AssumePrime = 1;
	end	else if (num==16'd14771) begin
		AssumePrime = 1;
	end	else if (num==16'd14779) begin
		AssumePrime = 1;
	end	else if (num==16'd14783) begin
		AssumePrime = 1;
	end	else if (num==16'd14797) begin
		AssumePrime = 1;
	end	else if (num==16'd14813) begin
		AssumePrime = 1;
	end	else if (num==16'd14821) begin
		AssumePrime = 1;
	end	else if (num==16'd14827) begin
		AssumePrime = 1;
	end	else if (num==16'd14831) begin
		AssumePrime = 1;
	end	else if (num==16'd14843) begin
		AssumePrime = 1;
	end	else if (num==16'd14851) begin
		AssumePrime = 1;
	end	else if (num==16'd14867) begin
		AssumePrime = 1;
	end	else if (num==16'd14869) begin
		AssumePrime = 1;
	end	else if (num==16'd14879) begin
		AssumePrime = 1;
	end	else if (num==16'd14887) begin
		AssumePrime = 1;
	end	else if (num==16'd14891) begin
		AssumePrime = 1;
	end	else if (num==16'd14897) begin
		AssumePrime = 1;
	end	else if (num==16'd14923) begin
		AssumePrime = 1;
	end	else if (num==16'd14929) begin
		AssumePrime = 1;
	end	else if (num==16'd14939) begin
		AssumePrime = 1;
	end	else if (num==16'd14947) begin
		AssumePrime = 1;
	end	else if (num==16'd14951) begin
		AssumePrime = 1;
	end	else if (num==16'd14957) begin
		AssumePrime = 1;
	end	else if (num==16'd14969) begin
		AssumePrime = 1;
	end	else if (num==16'd14983) begin
		AssumePrime = 1;
	end	else if (num==16'd15013) begin
		AssumePrime = 1;
	end	else if (num==16'd15017) begin
		AssumePrime = 1;
	end	else if (num==16'd15031) begin
		AssumePrime = 1;
	end	else if (num==16'd15053) begin
		AssumePrime = 1;
	end	else if (num==16'd15061) begin
		AssumePrime = 1;
	end	else if (num==16'd15073) begin
		AssumePrime = 1;
	end	else if (num==16'd15077) begin
		AssumePrime = 1;
	end	else if (num==16'd15083) begin
		AssumePrime = 1;
	end	else if (num==16'd15091) begin
		AssumePrime = 1;
	end	else if (num==16'd15101) begin
		AssumePrime = 1;
	end	else if (num==16'd15107) begin
		AssumePrime = 1;
	end	else if (num==16'd15121) begin
		AssumePrime = 1;
	end	else if (num==16'd15131) begin
		AssumePrime = 1;
	end	else if (num==16'd15137) begin
		AssumePrime = 1;
	end	else if (num==16'd15139) begin
		AssumePrime = 1;
	end	else if (num==16'd15149) begin
		AssumePrime = 1;
	end	else if (num==16'd15161) begin
		AssumePrime = 1;
	end	else if (num==16'd15173) begin
		AssumePrime = 1;
	end	else if (num==16'd15187) begin
		AssumePrime = 1;
	end	else if (num==16'd15193) begin
		AssumePrime = 1;
	end	else if (num==16'd15199) begin
		AssumePrime = 1;
	end	else if (num==16'd15217) begin
		AssumePrime = 1;
	end	else if (num==16'd15227) begin
		AssumePrime = 1;
	end	else if (num==16'd15233) begin
		AssumePrime = 1;
	end	else if (num==16'd15241) begin
		AssumePrime = 1;
	end	else if (num==16'd15259) begin
		AssumePrime = 1;
	end	else if (num==16'd15263) begin
		AssumePrime = 1;
	end	else if (num==16'd15269) begin
		AssumePrime = 1;
	end	else if (num==16'd15271) begin
		AssumePrime = 1;
	end	else if (num==16'd15277) begin
		AssumePrime = 1;
	end	else if (num==16'd15287) begin
		AssumePrime = 1;
	end	else if (num==16'd15289) begin
		AssumePrime = 1;
	end	else if (num==16'd15299) begin
		AssumePrime = 1;
	end	else if (num==16'd15307) begin
		AssumePrime = 1;
	end	else if (num==16'd15313) begin
		AssumePrime = 1;
	end	else if (num==16'd15319) begin
		AssumePrime = 1;
	end	else if (num==16'd15329) begin
		AssumePrime = 1;
	end	else if (num==16'd15331) begin
		AssumePrime = 1;
	end	else if (num==16'd15349) begin
		AssumePrime = 1;
	end	else if (num==16'd15359) begin
		AssumePrime = 1;
	end	else if (num==16'd15361) begin
		AssumePrime = 1;
	end	else if (num==16'd15373) begin
		AssumePrime = 1;
	end	else if (num==16'd15377) begin
		AssumePrime = 1;
	end	else if (num==16'd15383) begin
		AssumePrime = 1;
	end	else if (num==16'd15391) begin
		AssumePrime = 1;
	end	else if (num==16'd15401) begin
		AssumePrime = 1;
	end	else if (num==16'd15413) begin
		AssumePrime = 1;
	end	else if (num==16'd15427) begin
		AssumePrime = 1;
	end	else if (num==16'd15439) begin
		AssumePrime = 1;
	end	else if (num==16'd15443) begin
		AssumePrime = 1;
	end	else if (num==16'd15451) begin
		AssumePrime = 1;
	end	else if (num==16'd15461) begin
		AssumePrime = 1;
	end	else if (num==16'd15467) begin
		AssumePrime = 1;
	end	else if (num==16'd15473) begin
		AssumePrime = 1;
	end	else if (num==16'd15493) begin
		AssumePrime = 1;
	end	else if (num==16'd15497) begin
		AssumePrime = 1;
	end	else if (num==16'd15511) begin
		AssumePrime = 1;
	end	else if (num==16'd15527) begin
		AssumePrime = 1;
	end	else if (num==16'd15541) begin
		AssumePrime = 1;
	end	else if (num==16'd15551) begin
		AssumePrime = 1;
	end	else if (num==16'd15559) begin
		AssumePrime = 1;
	end	else if (num==16'd15569) begin
		AssumePrime = 1;
	end	else if (num==16'd15581) begin
		AssumePrime = 1;
	end	else if (num==16'd15583) begin
		AssumePrime = 1;
	end	else if (num==16'd15601) begin
		AssumePrime = 1;
	end	else if (num==16'd15607) begin
		AssumePrime = 1;
	end	else if (num==16'd15619) begin
		AssumePrime = 1;
	end	else if (num==16'd15629) begin
		AssumePrime = 1;
	end	else if (num==16'd15641) begin
		AssumePrime = 1;
	end	else if (num==16'd15643) begin
		AssumePrime = 1;
	end	else if (num==16'd15647) begin
		AssumePrime = 1;
	end	else if (num==16'd15649) begin
		AssumePrime = 1;
	end	else if (num==16'd15661) begin
		AssumePrime = 1;
	end	else if (num==16'd15667) begin
		AssumePrime = 1;
	end	else if (num==16'd15671) begin
		AssumePrime = 1;
	end	else if (num==16'd15679) begin
		AssumePrime = 1;
	end	else if (num==16'd15683) begin
		AssumePrime = 1;
	end	else if (num==16'd15727) begin
		AssumePrime = 1;
	end	else if (num==16'd15731) begin
		AssumePrime = 1;
	end	else if (num==16'd15733) begin
		AssumePrime = 1;
	end	else if (num==16'd15737) begin
		AssumePrime = 1;
	end	else if (num==16'd15739) begin
		AssumePrime = 1;
	end	else if (num==16'd15749) begin
		AssumePrime = 1;
	end	else if (num==16'd15761) begin
		AssumePrime = 1;
	end	else if (num==16'd15767) begin
		AssumePrime = 1;
	end	else if (num==16'd15773) begin
		AssumePrime = 1;
	end	else if (num==16'd15787) begin
		AssumePrime = 1;
	end	else if (num==16'd15791) begin
		AssumePrime = 1;
	end	else if (num==16'd15797) begin
		AssumePrime = 1;
	end	else if (num==16'd15803) begin
		AssumePrime = 1;
	end	else if (num==16'd15809) begin
		AssumePrime = 1;
	end	else if (num==16'd15817) begin
		AssumePrime = 1;
	end	else if (num==16'd15823) begin
		AssumePrime = 1;
	end	else if (num==16'd15859) begin
		AssumePrime = 1;
	end	else if (num==16'd15877) begin
		AssumePrime = 1;
	end	else if (num==16'd15881) begin
		AssumePrime = 1;
	end	else if (num==16'd15887) begin
		AssumePrime = 1;
	end	else if (num==16'd15889) begin
		AssumePrime = 1;
	end	else if (num==16'd15901) begin
		AssumePrime = 1;
	end	else if (num==16'd15907) begin
		AssumePrime = 1;
	end	else if (num==16'd15913) begin
		AssumePrime = 1;
	end	else if (num==16'd15919) begin
		AssumePrime = 1;
	end	else if (num==16'd15923) begin
		AssumePrime = 1;
	end	else if (num==16'd15937) begin
		AssumePrime = 1;
	end	else if (num==16'd15959) begin
		AssumePrime = 1;
	end	else if (num==16'd15971) begin
		AssumePrime = 1;
	end	else if (num==16'd15973) begin
		AssumePrime = 1;
	end	else if (num==16'd15991) begin
		AssumePrime = 1;
	end	else if (num==16'd16001) begin
		AssumePrime = 1;
	end	else if (num==16'd16007) begin
		AssumePrime = 1;
	end	else if (num==16'd16033) begin
		AssumePrime = 1;
	end	else if (num==16'd16057) begin
		AssumePrime = 1;
	end	else if (num==16'd16061) begin
		AssumePrime = 1;
	end	else if (num==16'd16063) begin
		AssumePrime = 1;
	end	else if (num==16'd16067) begin
		AssumePrime = 1;
	end	else if (num==16'd16069) begin
		AssumePrime = 1;
	end	else if (num==16'd16073) begin
		AssumePrime = 1;
	end	else if (num==16'd16087) begin
		AssumePrime = 1;
	end	else if (num==16'd16091) begin
		AssumePrime = 1;
	end	else if (num==16'd16097) begin
		AssumePrime = 1;
	end	else if (num==16'd16103) begin
		AssumePrime = 1;
	end	else if (num==16'd16111) begin
		AssumePrime = 1;
	end	else if (num==16'd16127) begin
		AssumePrime = 1;
	end	else if (num==16'd16139) begin
		AssumePrime = 1;
	end	else if (num==16'd16141) begin
		AssumePrime = 1;
	end	else if (num==16'd16183) begin
		AssumePrime = 1;
	end	else if (num==16'd16187) begin
		AssumePrime = 1;
	end	else if (num==16'd16189) begin
		AssumePrime = 1;
	end	else if (num==16'd16193) begin
		AssumePrime = 1;
	end	else if (num==16'd16217) begin
		AssumePrime = 1;
	end	else if (num==16'd16223) begin
		AssumePrime = 1;
	end	else if (num==16'd16229) begin
		AssumePrime = 1;
	end	else if (num==16'd16231) begin
		AssumePrime = 1;
	end	else if (num==16'd16249) begin
		AssumePrime = 1;
	end	else if (num==16'd16253) begin
		AssumePrime = 1;
	end	else if (num==16'd16267) begin
		AssumePrime = 1;
	end	else if (num==16'd16273) begin
		AssumePrime = 1;
	end	else if (num==16'd16301) begin
		AssumePrime = 1;
	end	else if (num==16'd16319) begin
		AssumePrime = 1;
	end	else if (num==16'd16333) begin
		AssumePrime = 1;
	end	else if (num==16'd16339) begin
		AssumePrime = 1;
	end	else if (num==16'd16349) begin
		AssumePrime = 1;
	end	else if (num==16'd16361) begin
		AssumePrime = 1;
	end	else if (num==16'd16363) begin
		AssumePrime = 1;
	end	else if (num==16'd16369) begin
		AssumePrime = 1;
	end	else if (num==16'd16381) begin
		AssumePrime = 1;
	end	else if (num==16'd16411) begin
		AssumePrime = 1;
	end	else if (num==16'd16417) begin
		AssumePrime = 1;
	end	else if (num==16'd16421) begin
		AssumePrime = 1;
	end	else if (num==16'd16427) begin
		AssumePrime = 1;
	end	else if (num==16'd16433) begin
		AssumePrime = 1;
	end	else if (num==16'd16447) begin
		AssumePrime = 1;
	end	else if (num==16'd16451) begin
		AssumePrime = 1;
	end	else if (num==16'd16453) begin
		AssumePrime = 1;
	end	else if (num==16'd16477) begin
		AssumePrime = 1;
	end	else if (num==16'd16481) begin
		AssumePrime = 1;
	end	else if (num==16'd16487) begin
		AssumePrime = 1;
	end	else if (num==16'd16493) begin
		AssumePrime = 1;
	end	else if (num==16'd16519) begin
		AssumePrime = 1;
	end	else if (num==16'd16529) begin
		AssumePrime = 1;
	end	else if (num==16'd16547) begin
		AssumePrime = 1;
	end	else if (num==16'd16553) begin
		AssumePrime = 1;
	end	else if (num==16'd16561) begin
		AssumePrime = 1;
	end	else if (num==16'd16567) begin
		AssumePrime = 1;
	end	else if (num==16'd16573) begin
		AssumePrime = 1;
	end	else if (num==16'd16603) begin
		AssumePrime = 1;
	end	else if (num==16'd16607) begin
		AssumePrime = 1;
	end	else if (num==16'd16619) begin
		AssumePrime = 1;
	end	else if (num==16'd16631) begin
		AssumePrime = 1;
	end	else if (num==16'd16633) begin
		AssumePrime = 1;
	end	else if (num==16'd16649) begin
		AssumePrime = 1;
	end	else if (num==16'd16651) begin
		AssumePrime = 1;
	end	else if (num==16'd16657) begin
		AssumePrime = 1;
	end	else if (num==16'd16661) begin
		AssumePrime = 1;
	end	else if (num==16'd16673) begin
		AssumePrime = 1;
	end	else if (num==16'd16691) begin
		AssumePrime = 1;
	end	else if (num==16'd16693) begin
		AssumePrime = 1;
	end	else if (num==16'd16699) begin
		AssumePrime = 1;
	end	else if (num==16'd16703) begin
		AssumePrime = 1;
	end	else if (num==16'd16729) begin
		AssumePrime = 1;
	end	else if (num==16'd16741) begin
		AssumePrime = 1;
	end	else if (num==16'd16747) begin
		AssumePrime = 1;
	end	else if (num==16'd16759) begin
		AssumePrime = 1;
	end	else if (num==16'd16763) begin
		AssumePrime = 1;
	end	else if (num==16'd16787) begin
		AssumePrime = 1;
	end	else if (num==16'd16811) begin
		AssumePrime = 1;
	end	else if (num==16'd16823) begin
		AssumePrime = 1;
	end	else if (num==16'd16829) begin
		AssumePrime = 1;
	end	else if (num==16'd16831) begin
		AssumePrime = 1;
	end	else if (num==16'd16843) begin
		AssumePrime = 1;
	end	else if (num==16'd16871) begin
		AssumePrime = 1;
	end	else if (num==16'd16879) begin
		AssumePrime = 1;
	end	else if (num==16'd16883) begin
		AssumePrime = 1;
	end	else if (num==16'd16889) begin
		AssumePrime = 1;
	end	else if (num==16'd16901) begin
		AssumePrime = 1;
	end	else if (num==16'd16903) begin
		AssumePrime = 1;
	end	else if (num==16'd16921) begin
		AssumePrime = 1;
	end	else if (num==16'd16927) begin
		AssumePrime = 1;
	end	else if (num==16'd16931) begin
		AssumePrime = 1;
	end	else if (num==16'd16937) begin
		AssumePrime = 1;
	end	else if (num==16'd16943) begin
		AssumePrime = 1;
	end	else if (num==16'd16963) begin
		AssumePrime = 1;
	end	else if (num==16'd16979) begin
		AssumePrime = 1;
	end	else if (num==16'd16981) begin
		AssumePrime = 1;
	end	else if (num==16'd16987) begin
		AssumePrime = 1;
	end	else if (num==16'd16993) begin
		AssumePrime = 1;
	end	else if (num==16'd17011) begin
		AssumePrime = 1;
	end	else if (num==16'd17021) begin
		AssumePrime = 1;
	end	else if (num==16'd17027) begin
		AssumePrime = 1;
	end	else if (num==16'd17029) begin
		AssumePrime = 1;
	end	else if (num==16'd17033) begin
		AssumePrime = 1;
	end	else if (num==16'd17041) begin
		AssumePrime = 1;
	end	else if (num==16'd17047) begin
		AssumePrime = 1;
	end	else if (num==16'd17053) begin
		AssumePrime = 1;
	end	else if (num==16'd17077) begin
		AssumePrime = 1;
	end	else if (num==16'd17093) begin
		AssumePrime = 1;
	end	else if (num==16'd17099) begin
		AssumePrime = 1;
	end	else if (num==16'd17107) begin
		AssumePrime = 1;
	end	else if (num==16'd17117) begin
		AssumePrime = 1;
	end	else if (num==16'd17123) begin
		AssumePrime = 1;
	end	else if (num==16'd17137) begin
		AssumePrime = 1;
	end	else if (num==16'd17159) begin
		AssumePrime = 1;
	end	else if (num==16'd17167) begin
		AssumePrime = 1;
	end	else if (num==16'd17183) begin
		AssumePrime = 1;
	end	else if (num==16'd17189) begin
		AssumePrime = 1;
	end	else if (num==16'd17191) begin
		AssumePrime = 1;
	end	else if (num==16'd17203) begin
		AssumePrime = 1;
	end	else if (num==16'd17207) begin
		AssumePrime = 1;
	end	else if (num==16'd17209) begin
		AssumePrime = 1;
	end	else if (num==16'd17231) begin
		AssumePrime = 1;
	end	else if (num==16'd17239) begin
		AssumePrime = 1;
	end	else if (num==16'd17257) begin
		AssumePrime = 1;
	end	else if (num==16'd17291) begin
		AssumePrime = 1;
	end	else if (num==16'd17293) begin
		AssumePrime = 1;
	end	else if (num==16'd17299) begin
		AssumePrime = 1;
	end	else if (num==16'd17317) begin
		AssumePrime = 1;
	end	else if (num==16'd17321) begin
		AssumePrime = 1;
	end	else if (num==16'd17327) begin
		AssumePrime = 1;
	end	else if (num==16'd17333) begin
		AssumePrime = 1;
	end	else if (num==16'd17341) begin
		AssumePrime = 1;
	end	else if (num==16'd17351) begin
		AssumePrime = 1;
	end	else if (num==16'd17359) begin
		AssumePrime = 1;
	end	else if (num==16'd17377) begin
		AssumePrime = 1;
	end	else if (num==16'd17383) begin
		AssumePrime = 1;
	end	else if (num==16'd17387) begin
		AssumePrime = 1;
	end	else if (num==16'd17389) begin
		AssumePrime = 1;
	end	else if (num==16'd17393) begin
		AssumePrime = 1;
	end	else if (num==16'd17401) begin
		AssumePrime = 1;
	end	else if (num==16'd17417) begin
		AssumePrime = 1;
	end	else if (num==16'd17419) begin
		AssumePrime = 1;
	end	else if (num==16'd17431) begin
		AssumePrime = 1;
	end	else if (num==16'd17443) begin
		AssumePrime = 1;
	end	else if (num==16'd17449) begin
		AssumePrime = 1;
	end	else if (num==16'd17467) begin
		AssumePrime = 1;
	end	else if (num==16'd17471) begin
		AssumePrime = 1;
	end	else if (num==16'd17477) begin
		AssumePrime = 1;
	end	else if (num==16'd17483) begin
		AssumePrime = 1;
	end	else if (num==16'd17489) begin
		AssumePrime = 1;
	end	else if (num==16'd17491) begin
		AssumePrime = 1;
	end	else if (num==16'd17497) begin
		AssumePrime = 1;
	end	else if (num==16'd17509) begin
		AssumePrime = 1;
	end	else if (num==16'd17519) begin
		AssumePrime = 1;
	end	else if (num==16'd17539) begin
		AssumePrime = 1;
	end	else if (num==16'd17551) begin
		AssumePrime = 1;
	end	else if (num==16'd17569) begin
		AssumePrime = 1;
	end	else if (num==16'd17573) begin
		AssumePrime = 1;
	end	else if (num==16'd17579) begin
		AssumePrime = 1;
	end	else if (num==16'd17581) begin
		AssumePrime = 1;
	end	else if (num==16'd17597) begin
		AssumePrime = 1;
	end	else if (num==16'd17599) begin
		AssumePrime = 1;
	end	else if (num==16'd17609) begin
		AssumePrime = 1;
	end	else if (num==16'd17623) begin
		AssumePrime = 1;
	end	else if (num==16'd17627) begin
		AssumePrime = 1;
	end	else if (num==16'd17657) begin
		AssumePrime = 1;
	end	else if (num==16'd17659) begin
		AssumePrime = 1;
	end	else if (num==16'd17669) begin
		AssumePrime = 1;
	end	else if (num==16'd17681) begin
		AssumePrime = 1;
	end	else if (num==16'd17683) begin
		AssumePrime = 1;
	end	else if (num==16'd17707) begin
		AssumePrime = 1;
	end	else if (num==16'd17713) begin
		AssumePrime = 1;
	end	else if (num==16'd17729) begin
		AssumePrime = 1;
	end	else if (num==16'd17737) begin
		AssumePrime = 1;
	end	else if (num==16'd17747) begin
		AssumePrime = 1;
	end	else if (num==16'd17749) begin
		AssumePrime = 1;
	end	else if (num==16'd17761) begin
		AssumePrime = 1;
	end	else if (num==16'd17783) begin
		AssumePrime = 1;
	end	else if (num==16'd17789) begin
		AssumePrime = 1;
	end	else if (num==16'd17791) begin
		AssumePrime = 1;
	end	else if (num==16'd17807) begin
		AssumePrime = 1;
	end	else if (num==16'd17827) begin
		AssumePrime = 1;
	end	else if (num==16'd17837) begin
		AssumePrime = 1;
	end	else if (num==16'd17839) begin
		AssumePrime = 1;
	end	else if (num==16'd17851) begin
		AssumePrime = 1;
	end	else if (num==16'd17863) begin
		AssumePrime = 1;
	end	else if (num==16'd17881) begin
		AssumePrime = 1;
	end	else if (num==16'd17891) begin
		AssumePrime = 1;
	end	else if (num==16'd17903) begin
		AssumePrime = 1;
	end	else if (num==16'd17909) begin
		AssumePrime = 1;
	end	else if (num==16'd17911) begin
		AssumePrime = 1;
	end	else if (num==16'd17921) begin
		AssumePrime = 1;
	end	else if (num==16'd17923) begin
		AssumePrime = 1;
	end	else if (num==16'd17929) begin
		AssumePrime = 1;
	end	else if (num==16'd17939) begin
		AssumePrime = 1;
	end	else if (num==16'd17957) begin
		AssumePrime = 1;
	end	else if (num==16'd17959) begin
		AssumePrime = 1;
	end	else if (num==16'd17971) begin
		AssumePrime = 1;
	end	else if (num==16'd17977) begin
		AssumePrime = 1;
	end	else if (num==16'd17981) begin
		AssumePrime = 1;
	end	else if (num==16'd17987) begin
		AssumePrime = 1;
	end	else if (num==16'd17989) begin
		AssumePrime = 1;
	end	else if (num==16'd18013) begin
		AssumePrime = 1;
	end	else if (num==16'd18041) begin
		AssumePrime = 1;
	end	else if (num==16'd18043) begin
		AssumePrime = 1;
	end	else if (num==16'd18047) begin
		AssumePrime = 1;
	end	else if (num==16'd18049) begin
		AssumePrime = 1;
	end	else if (num==16'd18059) begin
		AssumePrime = 1;
	end	else if (num==16'd18061) begin
		AssumePrime = 1;
	end	else if (num==16'd18077) begin
		AssumePrime = 1;
	end	else if (num==16'd18089) begin
		AssumePrime = 1;
	end	else if (num==16'd18097) begin
		AssumePrime = 1;
	end	else if (num==16'd18119) begin
		AssumePrime = 1;
	end	else if (num==16'd18121) begin
		AssumePrime = 1;
	end	else if (num==16'd18127) begin
		AssumePrime = 1;
	end	else if (num==16'd18131) begin
		AssumePrime = 1;
	end	else if (num==16'd18133) begin
		AssumePrime = 1;
	end	else if (num==16'd18143) begin
		AssumePrime = 1;
	end	else if (num==16'd18149) begin
		AssumePrime = 1;
	end	else if (num==16'd18169) begin
		AssumePrime = 1;
	end	else if (num==16'd18181) begin
		AssumePrime = 1;
	end	else if (num==16'd18191) begin
		AssumePrime = 1;
	end	else if (num==16'd18199) begin
		AssumePrime = 1;
	end	else if (num==16'd18211) begin
		AssumePrime = 1;
	end	else if (num==16'd18217) begin
		AssumePrime = 1;
	end	else if (num==16'd18223) begin
		AssumePrime = 1;
	end	else if (num==16'd18229) begin
		AssumePrime = 1;
	end	else if (num==16'd18233) begin
		AssumePrime = 1;
	end	else if (num==16'd18251) begin
		AssumePrime = 1;
	end	else if (num==16'd18253) begin
		AssumePrime = 1;
	end	else if (num==16'd18257) begin
		AssumePrime = 1;
	end	else if (num==16'd18269) begin
		AssumePrime = 1;
	end	else if (num==16'd18287) begin
		AssumePrime = 1;
	end	else if (num==16'd18289) begin
		AssumePrime = 1;
	end	else if (num==16'd18301) begin
		AssumePrime = 1;
	end	else if (num==16'd18307) begin
		AssumePrime = 1;
	end	else if (num==16'd18311) begin
		AssumePrime = 1;
	end	else if (num==16'd18313) begin
		AssumePrime = 1;
	end	else if (num==16'd18329) begin
		AssumePrime = 1;
	end	else if (num==16'd18341) begin
		AssumePrime = 1;
	end	else if (num==16'd18353) begin
		AssumePrime = 1;
	end	else if (num==16'd18367) begin
		AssumePrime = 1;
	end	else if (num==16'd18371) begin
		AssumePrime = 1;
	end	else if (num==16'd18379) begin
		AssumePrime = 1;
	end	else if (num==16'd18397) begin
		AssumePrime = 1;
	end	else if (num==16'd18401) begin
		AssumePrime = 1;
	end	else if (num==16'd18413) begin
		AssumePrime = 1;
	end	else if (num==16'd18427) begin
		AssumePrime = 1;
	end	else if (num==16'd18433) begin
		AssumePrime = 1;
	end	else if (num==16'd18439) begin
		AssumePrime = 1;
	end	else if (num==16'd18443) begin
		AssumePrime = 1;
	end	else if (num==16'd18451) begin
		AssumePrime = 1;
	end	else if (num==16'd18457) begin
		AssumePrime = 1;
	end	else if (num==16'd18461) begin
		AssumePrime = 1;
	end	else if (num==16'd18481) begin
		AssumePrime = 1;
	end	else if (num==16'd18493) begin
		AssumePrime = 1;
	end	else if (num==16'd18503) begin
		AssumePrime = 1;
	end	else if (num==16'd18517) begin
		AssumePrime = 1;
	end	else if (num==16'd18521) begin
		AssumePrime = 1;
	end	else if (num==16'd18523) begin
		AssumePrime = 1;
	end	else if (num==16'd18539) begin
		AssumePrime = 1;
	end	else if (num==16'd18541) begin
		AssumePrime = 1;
	end	else if (num==16'd18553) begin
		AssumePrime = 1;
	end	else if (num==16'd18583) begin
		AssumePrime = 1;
	end	else if (num==16'd18587) begin
		AssumePrime = 1;
	end	else if (num==16'd18593) begin
		AssumePrime = 1;
	end	else if (num==16'd18617) begin
		AssumePrime = 1;
	end	else if (num==16'd18637) begin
		AssumePrime = 1;
	end	else if (num==16'd18661) begin
		AssumePrime = 1;
	end	else if (num==16'd18671) begin
		AssumePrime = 1;
	end	else if (num==16'd18679) begin
		AssumePrime = 1;
	end	else if (num==16'd18691) begin
		AssumePrime = 1;
	end	else if (num==16'd18701) begin
		AssumePrime = 1;
	end	else if (num==16'd18713) begin
		AssumePrime = 1;
	end	else if (num==16'd18719) begin
		AssumePrime = 1;
	end	else if (num==16'd18731) begin
		AssumePrime = 1;
	end	else if (num==16'd18743) begin
		AssumePrime = 1;
	end	else if (num==16'd18749) begin
		AssumePrime = 1;
	end	else if (num==16'd18757) begin
		AssumePrime = 1;
	end	else if (num==16'd18773) begin
		AssumePrime = 1;
	end	else if (num==16'd18787) begin
		AssumePrime = 1;
	end	else if (num==16'd18793) begin
		AssumePrime = 1;
	end	else if (num==16'd18797) begin
		AssumePrime = 1;
	end	else if (num==16'd18803) begin
		AssumePrime = 1;
	end	else if (num==16'd18839) begin
		AssumePrime = 1;
	end	else if (num==16'd18859) begin
		AssumePrime = 1;
	end	else if (num==16'd18869) begin
		AssumePrime = 1;
	end	else if (num==16'd18899) begin
		AssumePrime = 1;
	end	else if (num==16'd18911) begin
		AssumePrime = 1;
	end	else if (num==16'd18913) begin
		AssumePrime = 1;
	end	else if (num==16'd18917) begin
		AssumePrime = 1;
	end	else if (num==16'd18919) begin
		AssumePrime = 1;
	end	else if (num==16'd18947) begin
		AssumePrime = 1;
	end	else if (num==16'd18959) begin
		AssumePrime = 1;
	end	else if (num==16'd18973) begin
		AssumePrime = 1;
	end	else if (num==16'd18979) begin
		AssumePrime = 1;
	end	else if (num==16'd19001) begin
		AssumePrime = 1;
	end	else if (num==16'd19009) begin
		AssumePrime = 1;
	end	else if (num==16'd19013) begin
		AssumePrime = 1;
	end	else if (num==16'd19031) begin
		AssumePrime = 1;
	end	else if (num==16'd19037) begin
		AssumePrime = 1;
	end	else if (num==16'd19051) begin
		AssumePrime = 1;
	end	else if (num==16'd19069) begin
		AssumePrime = 1;
	end	else if (num==16'd19073) begin
		AssumePrime = 1;
	end	else if (num==16'd19079) begin
		AssumePrime = 1;
	end	else if (num==16'd19081) begin
		AssumePrime = 1;
	end	else if (num==16'd19087) begin
		AssumePrime = 1;
	end	else if (num==16'd19121) begin
		AssumePrime = 1;
	end	else if (num==16'd19139) begin
		AssumePrime = 1;
	end	else if (num==16'd19141) begin
		AssumePrime = 1;
	end	else if (num==16'd19157) begin
		AssumePrime = 1;
	end	else if (num==16'd19163) begin
		AssumePrime = 1;
	end	else if (num==16'd19181) begin
		AssumePrime = 1;
	end	else if (num==16'd19183) begin
		AssumePrime = 1;
	end	else if (num==16'd19207) begin
		AssumePrime = 1;
	end	else if (num==16'd19211) begin
		AssumePrime = 1;
	end	else if (num==16'd19213) begin
		AssumePrime = 1;
	end	else if (num==16'd19219) begin
		AssumePrime = 1;
	end	else if (num==16'd19231) begin
		AssumePrime = 1;
	end	else if (num==16'd19237) begin
		AssumePrime = 1;
	end	else if (num==16'd19249) begin
		AssumePrime = 1;
	end	else if (num==16'd19259) begin
		AssumePrime = 1;
	end	else if (num==16'd19267) begin
		AssumePrime = 1;
	end	else if (num==16'd19273) begin
		AssumePrime = 1;
	end	else if (num==16'd19289) begin
		AssumePrime = 1;
	end	else if (num==16'd19301) begin
		AssumePrime = 1;
	end	else if (num==16'd19309) begin
		AssumePrime = 1;
	end	else if (num==16'd19319) begin
		AssumePrime = 1;
	end	else if (num==16'd19333) begin
		AssumePrime = 1;
	end	else if (num==16'd19373) begin
		AssumePrime = 1;
	end	else if (num==16'd19379) begin
		AssumePrime = 1;
	end	else if (num==16'd19381) begin
		AssumePrime = 1;
	end	else if (num==16'd19387) begin
		AssumePrime = 1;
	end	else if (num==16'd19391) begin
		AssumePrime = 1;
	end	else if (num==16'd19403) begin
		AssumePrime = 1;
	end	else if (num==16'd19417) begin
		AssumePrime = 1;
	end	else if (num==16'd19421) begin
		AssumePrime = 1;
	end	else if (num==16'd19423) begin
		AssumePrime = 1;
	end	else if (num==16'd19427) begin
		AssumePrime = 1;
	end	else if (num==16'd19429) begin
		AssumePrime = 1;
	end	else if (num==16'd19433) begin
		AssumePrime = 1;
	end	else if (num==16'd19441) begin
		AssumePrime = 1;
	end	else if (num==16'd19447) begin
		AssumePrime = 1;
	end	else if (num==16'd19457) begin
		AssumePrime = 1;
	end	else if (num==16'd19463) begin
		AssumePrime = 1;
	end	else if (num==16'd19469) begin
		AssumePrime = 1;
	end	else if (num==16'd19471) begin
		AssumePrime = 1;
	end	else if (num==16'd19477) begin
		AssumePrime = 1;
	end	else if (num==16'd19483) begin
		AssumePrime = 1;
	end	else if (num==16'd19489) begin
		AssumePrime = 1;
	end	else if (num==16'd19501) begin
		AssumePrime = 1;
	end	else if (num==16'd19507) begin
		AssumePrime = 1;
	end	else if (num==16'd19531) begin
		AssumePrime = 1;
	end	else if (num==16'd19541) begin
		AssumePrime = 1;
	end	else if (num==16'd19543) begin
		AssumePrime = 1;
	end	else if (num==16'd19553) begin
		AssumePrime = 1;
	end	else if (num==16'd19559) begin
		AssumePrime = 1;
	end	else if (num==16'd19571) begin
		AssumePrime = 1;
	end	else if (num==16'd19577) begin
		AssumePrime = 1;
	end	else if (num==16'd19583) begin
		AssumePrime = 1;
	end	else if (num==16'd19597) begin
		AssumePrime = 1;
	end	else if (num==16'd19603) begin
		AssumePrime = 1;
	end	else if (num==16'd19609) begin
		AssumePrime = 1;
	end	else if (num==16'd19661) begin
		AssumePrime = 1;
	end	else if (num==16'd19681) begin
		AssumePrime = 1;
	end	else if (num==16'd19687) begin
		AssumePrime = 1;
	end	else if (num==16'd19697) begin
		AssumePrime = 1;
	end	else if (num==16'd19699) begin
		AssumePrime = 1;
	end	else if (num==16'd19709) begin
		AssumePrime = 1;
	end	else if (num==16'd19717) begin
		AssumePrime = 1;
	end	else if (num==16'd19727) begin
		AssumePrime = 1;
	end	else if (num==16'd19739) begin
		AssumePrime = 1;
	end	else if (num==16'd19751) begin
		AssumePrime = 1;
	end	else if (num==16'd19753) begin
		AssumePrime = 1;
	end	else if (num==16'd19759) begin
		AssumePrime = 1;
	end	else if (num==16'd19763) begin
		AssumePrime = 1;
	end	else if (num==16'd19777) begin
		AssumePrime = 1;
	end	else if (num==16'd19793) begin
		AssumePrime = 1;
	end	else if (num==16'd19801) begin
		AssumePrime = 1;
	end	else if (num==16'd19813) begin
		AssumePrime = 1;
	end	else if (num==16'd19819) begin
		AssumePrime = 1;
	end	else if (num==16'd19841) begin
		AssumePrime = 1;
	end	else if (num==16'd19843) begin
		AssumePrime = 1;
	end	else if (num==16'd19853) begin
		AssumePrime = 1;
	end	else if (num==16'd19861) begin
		AssumePrime = 1;
	end	else if (num==16'd19867) begin
		AssumePrime = 1;
	end	else if (num==16'd19889) begin
		AssumePrime = 1;
	end	else if (num==16'd19891) begin
		AssumePrime = 1;
	end	else if (num==16'd19913) begin
		AssumePrime = 1;
	end	else if (num==16'd19919) begin
		AssumePrime = 1;
	end	else if (num==16'd19927) begin
		AssumePrime = 1;
	end	else if (num==16'd19937) begin
		AssumePrime = 1;
	end	else if (num==16'd19949) begin
		AssumePrime = 1;
	end	else if (num==16'd19961) begin
		AssumePrime = 1;
	end	else if (num==16'd19963) begin
		AssumePrime = 1;
	end	else if (num==16'd19973) begin
		AssumePrime = 1;
	end	else if (num==16'd19979) begin
		AssumePrime = 1;
	end	else if (num==16'd19991) begin
		AssumePrime = 1;
	end	else if (num==16'd19993) begin
		AssumePrime = 1;
	end	else if (num==16'd19997) begin
		AssumePrime = 1;
	end	else if (num==16'd20011) begin
		AssumePrime = 1;
	end	else if (num==16'd20021) begin
		AssumePrime = 1;
	end	else if (num==16'd20023) begin
		AssumePrime = 1;
	end	else if (num==16'd20029) begin
		AssumePrime = 1;
	end	else if (num==16'd20047) begin
		AssumePrime = 1;
	end	else if (num==16'd20051) begin
		AssumePrime = 1;
	end	else if (num==16'd20063) begin
		AssumePrime = 1;
	end	else if (num==16'd20071) begin
		AssumePrime = 1;
	end	else if (num==16'd20089) begin
		AssumePrime = 1;
	end	else if (num==16'd20101) begin
		AssumePrime = 1;
	end	else if (num==16'd20107) begin
		AssumePrime = 1;
	end	else if (num==16'd20113) begin
		AssumePrime = 1;
	end	else if (num==16'd20117) begin
		AssumePrime = 1;
	end	else if (num==16'd20123) begin
		AssumePrime = 1;
	end	else if (num==16'd20129) begin
		AssumePrime = 1;
	end	else if (num==16'd20143) begin
		AssumePrime = 1;
	end	else if (num==16'd20147) begin
		AssumePrime = 1;
	end	else if (num==16'd20149) begin
		AssumePrime = 1;
	end	else if (num==16'd20161) begin
		AssumePrime = 1;
	end	else if (num==16'd20173) begin
		AssumePrime = 1;
	end	else if (num==16'd20177) begin
		AssumePrime = 1;
	end	else if (num==16'd20183) begin
		AssumePrime = 1;
	end	else if (num==16'd20201) begin
		AssumePrime = 1;
	end	else if (num==16'd20219) begin
		AssumePrime = 1;
	end	else if (num==16'd20231) begin
		AssumePrime = 1;
	end	else if (num==16'd20233) begin
		AssumePrime = 1;
	end	else if (num==16'd20249) begin
		AssumePrime = 1;
	end	else if (num==16'd20261) begin
		AssumePrime = 1;
	end	else if (num==16'd20269) begin
		AssumePrime = 1;
	end	else if (num==16'd20287) begin
		AssumePrime = 1;
	end	else if (num==16'd20297) begin
		AssumePrime = 1;
	end	else if (num==16'd20323) begin
		AssumePrime = 1;
	end	else if (num==16'd20327) begin
		AssumePrime = 1;
	end	else if (num==16'd20333) begin
		AssumePrime = 1;
	end	else if (num==16'd20341) begin
		AssumePrime = 1;
	end	else if (num==16'd20347) begin
		AssumePrime = 1;
	end	else if (num==16'd20353) begin
		AssumePrime = 1;
	end	else if (num==16'd20357) begin
		AssumePrime = 1;
	end	else if (num==16'd20359) begin
		AssumePrime = 1;
	end	else if (num==16'd20369) begin
		AssumePrime = 1;
	end	else if (num==16'd20389) begin
		AssumePrime = 1;
	end	else if (num==16'd20393) begin
		AssumePrime = 1;
	end	else if (num==16'd20399) begin
		AssumePrime = 1;
	end	else if (num==16'd20407) begin
		AssumePrime = 1;
	end	else if (num==16'd20411) begin
		AssumePrime = 1;
	end	else if (num==16'd20431) begin
		AssumePrime = 1;
	end	else if (num==16'd20441) begin
		AssumePrime = 1;
	end	else if (num==16'd20443) begin
		AssumePrime = 1;
	end	else if (num==16'd20477) begin
		AssumePrime = 1;
	end	else if (num==16'd20479) begin
		AssumePrime = 1;
	end	else if (num==16'd20483) begin
		AssumePrime = 1;
	end	else if (num==16'd20507) begin
		AssumePrime = 1;
	end	else if (num==16'd20509) begin
		AssumePrime = 1;
	end	else if (num==16'd20521) begin
		AssumePrime = 1;
	end	else if (num==16'd20533) begin
		AssumePrime = 1;
	end	else if (num==16'd20543) begin
		AssumePrime = 1;
	end	else if (num==16'd20549) begin
		AssumePrime = 1;
	end	else if (num==16'd20551) begin
		AssumePrime = 1;
	end	else if (num==16'd20563) begin
		AssumePrime = 1;
	end	else if (num==16'd20593) begin
		AssumePrime = 1;
	end	else if (num==16'd20599) begin
		AssumePrime = 1;
	end	else if (num==16'd20611) begin
		AssumePrime = 1;
	end	else if (num==16'd20627) begin
		AssumePrime = 1;
	end	else if (num==16'd20639) begin
		AssumePrime = 1;
	end	else if (num==16'd20641) begin
		AssumePrime = 1;
	end	else if (num==16'd20663) begin
		AssumePrime = 1;
	end	else if (num==16'd20681) begin
		AssumePrime = 1;
	end	else if (num==16'd20693) begin
		AssumePrime = 1;
	end	else if (num==16'd20707) begin
		AssumePrime = 1;
	end	else if (num==16'd20717) begin
		AssumePrime = 1;
	end	else if (num==16'd20719) begin
		AssumePrime = 1;
	end	else if (num==16'd20731) begin
		AssumePrime = 1;
	end	else if (num==16'd20743) begin
		AssumePrime = 1;
	end	else if (num==16'd20747) begin
		AssumePrime = 1;
	end	else if (num==16'd20749) begin
		AssumePrime = 1;
	end	else if (num==16'd20753) begin
		AssumePrime = 1;
	end	else if (num==16'd20759) begin
		AssumePrime = 1;
	end	else if (num==16'd20771) begin
		AssumePrime = 1;
	end	else if (num==16'd20773) begin
		AssumePrime = 1;
	end	else if (num==16'd20789) begin
		AssumePrime = 1;
	end	else if (num==16'd20807) begin
		AssumePrime = 1;
	end	else if (num==16'd20809) begin
		AssumePrime = 1;
	end	else if (num==16'd20849) begin
		AssumePrime = 1;
	end	else if (num==16'd20857) begin
		AssumePrime = 1;
	end	else if (num==16'd20873) begin
		AssumePrime = 1;
	end	else if (num==16'd20879) begin
		AssumePrime = 1;
	end	else if (num==16'd20887) begin
		AssumePrime = 1;
	end	else if (num==16'd20897) begin
		AssumePrime = 1;
	end	else if (num==16'd20899) begin
		AssumePrime = 1;
	end	else if (num==16'd20903) begin
		AssumePrime = 1;
	end	else if (num==16'd20921) begin
		AssumePrime = 1;
	end	else if (num==16'd20929) begin
		AssumePrime = 1;
	end	else if (num==16'd20939) begin
		AssumePrime = 1;
	end	else if (num==16'd20947) begin
		AssumePrime = 1;
	end	else if (num==16'd20959) begin
		AssumePrime = 1;
	end	else if (num==16'd20963) begin
		AssumePrime = 1;
	end	else if (num==16'd20981) begin
		AssumePrime = 1;
	end	else if (num==16'd20983) begin
		AssumePrime = 1;
	end	else if (num==16'd21001) begin
		AssumePrime = 1;
	end	else if (num==16'd21011) begin
		AssumePrime = 1;
	end	else if (num==16'd21013) begin
		AssumePrime = 1;
	end	else if (num==16'd21017) begin
		AssumePrime = 1;
	end	else if (num==16'd21019) begin
		AssumePrime = 1;
	end	else if (num==16'd21023) begin
		AssumePrime = 1;
	end	else if (num==16'd21031) begin
		AssumePrime = 1;
	end	else if (num==16'd21059) begin
		AssumePrime = 1;
	end	else if (num==16'd21061) begin
		AssumePrime = 1;
	end	else if (num==16'd21067) begin
		AssumePrime = 1;
	end	else if (num==16'd21089) begin
		AssumePrime = 1;
	end	else if (num==16'd21101) begin
		AssumePrime = 1;
	end	else if (num==16'd21107) begin
		AssumePrime = 1;
	end	else if (num==16'd21121) begin
		AssumePrime = 1;
	end	else if (num==16'd21139) begin
		AssumePrime = 1;
	end	else if (num==16'd21143) begin
		AssumePrime = 1;
	end	else if (num==16'd21149) begin
		AssumePrime = 1;
	end	else if (num==16'd21157) begin
		AssumePrime = 1;
	end	else if (num==16'd21163) begin
		AssumePrime = 1;
	end	else if (num==16'd21169) begin
		AssumePrime = 1;
	end	else if (num==16'd21179) begin
		AssumePrime = 1;
	end	else if (num==16'd21187) begin
		AssumePrime = 1;
	end	else if (num==16'd21191) begin
		AssumePrime = 1;
	end	else if (num==16'd21193) begin
		AssumePrime = 1;
	end	else if (num==16'd21211) begin
		AssumePrime = 1;
	end	else if (num==16'd21221) begin
		AssumePrime = 1;
	end	else if (num==16'd21227) begin
		AssumePrime = 1;
	end	else if (num==16'd21247) begin
		AssumePrime = 1;
	end	else if (num==16'd21269) begin
		AssumePrime = 1;
	end	else if (num==16'd21277) begin
		AssumePrime = 1;
	end	else if (num==16'd21283) begin
		AssumePrime = 1;
	end	else if (num==16'd21313) begin
		AssumePrime = 1;
	end	else if (num==16'd21317) begin
		AssumePrime = 1;
	end	else if (num==16'd21319) begin
		AssumePrime = 1;
	end	else if (num==16'd21323) begin
		AssumePrime = 1;
	end	else if (num==16'd21341) begin
		AssumePrime = 1;
	end	else if (num==16'd21347) begin
		AssumePrime = 1;
	end	else if (num==16'd21377) begin
		AssumePrime = 1;
	end	else if (num==16'd21379) begin
		AssumePrime = 1;
	end	else if (num==16'd21383) begin
		AssumePrime = 1;
	end	else if (num==16'd21391) begin
		AssumePrime = 1;
	end	else if (num==16'd21397) begin
		AssumePrime = 1;
	end	else if (num==16'd21401) begin
		AssumePrime = 1;
	end	else if (num==16'd21407) begin
		AssumePrime = 1;
	end	else if (num==16'd21419) begin
		AssumePrime = 1;
	end	else if (num==16'd21433) begin
		AssumePrime = 1;
	end	else if (num==16'd21467) begin
		AssumePrime = 1;
	end	else if (num==16'd21481) begin
		AssumePrime = 1;
	end	else if (num==16'd21487) begin
		AssumePrime = 1;
	end	else if (num==16'd21491) begin
		AssumePrime = 1;
	end	else if (num==16'd21493) begin
		AssumePrime = 1;
	end	else if (num==16'd21499) begin
		AssumePrime = 1;
	end	else if (num==16'd21503) begin
		AssumePrime = 1;
	end	else if (num==16'd21517) begin
		AssumePrime = 1;
	end	else if (num==16'd21521) begin
		AssumePrime = 1;
	end	else if (num==16'd21523) begin
		AssumePrime = 1;
	end	else if (num==16'd21529) begin
		AssumePrime = 1;
	end	else if (num==16'd21557) begin
		AssumePrime = 1;
	end	else if (num==16'd21559) begin
		AssumePrime = 1;
	end	else if (num==16'd21563) begin
		AssumePrime = 1;
	end	else if (num==16'd21569) begin
		AssumePrime = 1;
	end	else if (num==16'd21577) begin
		AssumePrime = 1;
	end	else if (num==16'd21587) begin
		AssumePrime = 1;
	end	else if (num==16'd21589) begin
		AssumePrime = 1;
	end	else if (num==16'd21599) begin
		AssumePrime = 1;
	end	else if (num==16'd21601) begin
		AssumePrime = 1;
	end	else if (num==16'd21611) begin
		AssumePrime = 1;
	end	else if (num==16'd21613) begin
		AssumePrime = 1;
	end	else if (num==16'd21617) begin
		AssumePrime = 1;
	end	else if (num==16'd21647) begin
		AssumePrime = 1;
	end	else if (num==16'd21649) begin
		AssumePrime = 1;
	end	else if (num==16'd21661) begin
		AssumePrime = 1;
	end	else if (num==16'd21673) begin
		AssumePrime = 1;
	end	else if (num==16'd21683) begin
		AssumePrime = 1;
	end	else if (num==16'd21701) begin
		AssumePrime = 1;
	end	else if (num==16'd21713) begin
		AssumePrime = 1;
	end	else if (num==16'd21727) begin
		AssumePrime = 1;
	end	else if (num==16'd21737) begin
		AssumePrime = 1;
	end	else if (num==16'd21739) begin
		AssumePrime = 1;
	end	else if (num==16'd21751) begin
		AssumePrime = 1;
	end	else if (num==16'd21757) begin
		AssumePrime = 1;
	end	else if (num==16'd21767) begin
		AssumePrime = 1;
	end	else if (num==16'd21773) begin
		AssumePrime = 1;
	end	else if (num==16'd21787) begin
		AssumePrime = 1;
	end	else if (num==16'd21799) begin
		AssumePrime = 1;
	end	else if (num==16'd21803) begin
		AssumePrime = 1;
	end	else if (num==16'd21817) begin
		AssumePrime = 1;
	end	else if (num==16'd21821) begin
		AssumePrime = 1;
	end	else if (num==16'd21839) begin
		AssumePrime = 1;
	end	else if (num==16'd21841) begin
		AssumePrime = 1;
	end	else if (num==16'd21851) begin
		AssumePrime = 1;
	end	else if (num==16'd21859) begin
		AssumePrime = 1;
	end	else if (num==16'd21863) begin
		AssumePrime = 1;
	end	else if (num==16'd21871) begin
		AssumePrime = 1;
	end	else if (num==16'd21881) begin
		AssumePrime = 1;
	end	else if (num==16'd21893) begin
		AssumePrime = 1;
	end	else if (num==16'd21911) begin
		AssumePrime = 1;
	end	else if (num==16'd21929) begin
		AssumePrime = 1;
	end	else if (num==16'd21937) begin
		AssumePrime = 1;
	end	else if (num==16'd21943) begin
		AssumePrime = 1;
	end	else if (num==16'd21961) begin
		AssumePrime = 1;
	end	else if (num==16'd21977) begin
		AssumePrime = 1;
	end	else if (num==16'd21991) begin
		AssumePrime = 1;
	end	else if (num==16'd21997) begin
		AssumePrime = 1;
	end	else if (num==16'd22003) begin
		AssumePrime = 1;
	end	else if (num==16'd22013) begin
		AssumePrime = 1;
	end	else if (num==16'd22027) begin
		AssumePrime = 1;
	end	else if (num==16'd22031) begin
		AssumePrime = 1;
	end	else if (num==16'd22037) begin
		AssumePrime = 1;
	end	else if (num==16'd22039) begin
		AssumePrime = 1;
	end	else if (num==16'd22051) begin
		AssumePrime = 1;
	end	else if (num==16'd22063) begin
		AssumePrime = 1;
	end	else if (num==16'd22067) begin
		AssumePrime = 1;
	end	else if (num==16'd22073) begin
		AssumePrime = 1;
	end	else if (num==16'd22079) begin
		AssumePrime = 1;
	end	else if (num==16'd22091) begin
		AssumePrime = 1;
	end	else if (num==16'd22093) begin
		AssumePrime = 1;
	end	else if (num==16'd22109) begin
		AssumePrime = 1;
	end	else if (num==16'd22111) begin
		AssumePrime = 1;
	end	else if (num==16'd22123) begin
		AssumePrime = 1;
	end	else if (num==16'd22129) begin
		AssumePrime = 1;
	end	else if (num==16'd22133) begin
		AssumePrime = 1;
	end	else if (num==16'd22147) begin
		AssumePrime = 1;
	end	else if (num==16'd22153) begin
		AssumePrime = 1;
	end	else if (num==16'd22157) begin
		AssumePrime = 1;
	end	else if (num==16'd22159) begin
		AssumePrime = 1;
	end	else if (num==16'd22171) begin
		AssumePrime = 1;
	end	else if (num==16'd22189) begin
		AssumePrime = 1;
	end	else if (num==16'd22193) begin
		AssumePrime = 1;
	end	else if (num==16'd22229) begin
		AssumePrime = 1;
	end	else if (num==16'd22247) begin
		AssumePrime = 1;
	end	else if (num==16'd22259) begin
		AssumePrime = 1;
	end	else if (num==16'd22271) begin
		AssumePrime = 1;
	end	else if (num==16'd22273) begin
		AssumePrime = 1;
	end	else if (num==16'd22277) begin
		AssumePrime = 1;
	end	else if (num==16'd22279) begin
		AssumePrime = 1;
	end	else if (num==16'd22283) begin
		AssumePrime = 1;
	end	else if (num==16'd22291) begin
		AssumePrime = 1;
	end	else if (num==16'd22303) begin
		AssumePrime = 1;
	end	else if (num==16'd22307) begin
		AssumePrime = 1;
	end	else if (num==16'd22343) begin
		AssumePrime = 1;
	end	else if (num==16'd22349) begin
		AssumePrime = 1;
	end	else if (num==16'd22367) begin
		AssumePrime = 1;
	end	else if (num==16'd22369) begin
		AssumePrime = 1;
	end	else if (num==16'd22381) begin
		AssumePrime = 1;
	end	else if (num==16'd22391) begin
		AssumePrime = 1;
	end	else if (num==16'd22397) begin
		AssumePrime = 1;
	end	else if (num==16'd22409) begin
		AssumePrime = 1;
	end	else if (num==16'd22433) begin
		AssumePrime = 1;
	end	else if (num==16'd22441) begin
		AssumePrime = 1;
	end	else if (num==16'd22447) begin
		AssumePrime = 1;
	end	else if (num==16'd22453) begin
		AssumePrime = 1;
	end	else if (num==16'd22469) begin
		AssumePrime = 1;
	end	else if (num==16'd22481) begin
		AssumePrime = 1;
	end	else if (num==16'd22483) begin
		AssumePrime = 1;
	end	else if (num==16'd22501) begin
		AssumePrime = 1;
	end	else if (num==16'd22511) begin
		AssumePrime = 1;
	end	else if (num==16'd22531) begin
		AssumePrime = 1;
	end	else if (num==16'd22541) begin
		AssumePrime = 1;
	end	else if (num==16'd22543) begin
		AssumePrime = 1;
	end	else if (num==16'd22549) begin
		AssumePrime = 1;
	end	else if (num==16'd22567) begin
		AssumePrime = 1;
	end	else if (num==16'd22571) begin
		AssumePrime = 1;
	end	else if (num==16'd22573) begin
		AssumePrime = 1;
	end	else if (num==16'd22613) begin
		AssumePrime = 1;
	end	else if (num==16'd22619) begin
		AssumePrime = 1;
	end	else if (num==16'd22621) begin
		AssumePrime = 1;
	end	else if (num==16'd22637) begin
		AssumePrime = 1;
	end	else if (num==16'd22639) begin
		AssumePrime = 1;
	end	else if (num==16'd22643) begin
		AssumePrime = 1;
	end	else if (num==16'd22651) begin
		AssumePrime = 1;
	end	else if (num==16'd22669) begin
		AssumePrime = 1;
	end	else if (num==16'd22679) begin
		AssumePrime = 1;
	end	else if (num==16'd22691) begin
		AssumePrime = 1;
	end	else if (num==16'd22697) begin
		AssumePrime = 1;
	end	else if (num==16'd22699) begin
		AssumePrime = 1;
	end	else if (num==16'd22709) begin
		AssumePrime = 1;
	end	else if (num==16'd22717) begin
		AssumePrime = 1;
	end	else if (num==16'd22721) begin
		AssumePrime = 1;
	end	else if (num==16'd22727) begin
		AssumePrime = 1;
	end	else if (num==16'd22739) begin
		AssumePrime = 1;
	end	else if (num==16'd22741) begin
		AssumePrime = 1;
	end	else if (num==16'd22751) begin
		AssumePrime = 1;
	end	else if (num==16'd22769) begin
		AssumePrime = 1;
	end	else if (num==16'd22777) begin
		AssumePrime = 1;
	end	else if (num==16'd22783) begin
		AssumePrime = 1;
	end	else if (num==16'd22787) begin
		AssumePrime = 1;
	end	else if (num==16'd22807) begin
		AssumePrime = 1;
	end	else if (num==16'd22811) begin
		AssumePrime = 1;
	end	else if (num==16'd22817) begin
		AssumePrime = 1;
	end	else if (num==16'd22853) begin
		AssumePrime = 1;
	end	else if (num==16'd22859) begin
		AssumePrime = 1;
	end	else if (num==16'd22861) begin
		AssumePrime = 1;
	end	else if (num==16'd22871) begin
		AssumePrime = 1;
	end	else if (num==16'd22877) begin
		AssumePrime = 1;
	end	else if (num==16'd22901) begin
		AssumePrime = 1;
	end	else if (num==16'd22907) begin
		AssumePrime = 1;
	end	else if (num==16'd22921) begin
		AssumePrime = 1;
	end	else if (num==16'd22937) begin
		AssumePrime = 1;
	end	else if (num==16'd22943) begin
		AssumePrime = 1;
	end	else if (num==16'd22961) begin
		AssumePrime = 1;
	end	else if (num==16'd22963) begin
		AssumePrime = 1;
	end	else if (num==16'd22973) begin
		AssumePrime = 1;
	end	else if (num==16'd22993) begin
		AssumePrime = 1;
	end	else if (num==16'd23003) begin
		AssumePrime = 1;
	end	else if (num==16'd23011) begin
		AssumePrime = 1;
	end	else if (num==16'd23017) begin
		AssumePrime = 1;
	end	else if (num==16'd23021) begin
		AssumePrime = 1;
	end	else if (num==16'd23027) begin
		AssumePrime = 1;
	end	else if (num==16'd23029) begin
		AssumePrime = 1;
	end	else if (num==16'd23039) begin
		AssumePrime = 1;
	end	else if (num==16'd23041) begin
		AssumePrime = 1;
	end	else if (num==16'd23053) begin
		AssumePrime = 1;
	end	else if (num==16'd23057) begin
		AssumePrime = 1;
	end	else if (num==16'd23059) begin
		AssumePrime = 1;
	end	else if (num==16'd23063) begin
		AssumePrime = 1;
	end	else if (num==16'd23071) begin
		AssumePrime = 1;
	end	else if (num==16'd23081) begin
		AssumePrime = 1;
	end	else if (num==16'd23087) begin
		AssumePrime = 1;
	end	else if (num==16'd23099) begin
		AssumePrime = 1;
	end	else if (num==16'd23117) begin
		AssumePrime = 1;
	end	else if (num==16'd23131) begin
		AssumePrime = 1;
	end	else if (num==16'd23143) begin
		AssumePrime = 1;
	end	else if (num==16'd23159) begin
		AssumePrime = 1;
	end	else if (num==16'd23167) begin
		AssumePrime = 1;
	end	else if (num==16'd23173) begin
		AssumePrime = 1;
	end	else if (num==16'd23189) begin
		AssumePrime = 1;
	end	else if (num==16'd23197) begin
		AssumePrime = 1;
	end	else if (num==16'd23201) begin
		AssumePrime = 1;
	end	else if (num==16'd23203) begin
		AssumePrime = 1;
	end	else if (num==16'd23209) begin
		AssumePrime = 1;
	end	else if (num==16'd23227) begin
		AssumePrime = 1;
	end	else if (num==16'd23251) begin
		AssumePrime = 1;
	end	else if (num==16'd23269) begin
		AssumePrime = 1;
	end	else if (num==16'd23279) begin
		AssumePrime = 1;
	end	else if (num==16'd23291) begin
		AssumePrime = 1;
	end	else if (num==16'd23293) begin
		AssumePrime = 1;
	end	else if (num==16'd23297) begin
		AssumePrime = 1;
	end	else if (num==16'd23311) begin
		AssumePrime = 1;
	end	else if (num==16'd23321) begin
		AssumePrime = 1;
	end	else if (num==16'd23327) begin
		AssumePrime = 1;
	end	else if (num==16'd23333) begin
		AssumePrime = 1;
	end	else if (num==16'd23339) begin
		AssumePrime = 1;
	end	else if (num==16'd23357) begin
		AssumePrime = 1;
	end	else if (num==16'd23369) begin
		AssumePrime = 1;
	end	else if (num==16'd23371) begin
		AssumePrime = 1;
	end	else if (num==16'd23399) begin
		AssumePrime = 1;
	end	else if (num==16'd23417) begin
		AssumePrime = 1;
	end	else if (num==16'd23431) begin
		AssumePrime = 1;
	end	else if (num==16'd23447) begin
		AssumePrime = 1;
	end	else if (num==16'd23459) begin
		AssumePrime = 1;
	end	else if (num==16'd23473) begin
		AssumePrime = 1;
	end	else if (num==16'd23497) begin
		AssumePrime = 1;
	end	else if (num==16'd23509) begin
		AssumePrime = 1;
	end	else if (num==16'd23531) begin
		AssumePrime = 1;
	end	else if (num==16'd23537) begin
		AssumePrime = 1;
	end	else if (num==16'd23539) begin
		AssumePrime = 1;
	end	else if (num==16'd23549) begin
		AssumePrime = 1;
	end	else if (num==16'd23557) begin
		AssumePrime = 1;
	end	else if (num==16'd23561) begin
		AssumePrime = 1;
	end	else if (num==16'd23563) begin
		AssumePrime = 1;
	end	else if (num==16'd23567) begin
		AssumePrime = 1;
	end	else if (num==16'd23581) begin
		AssumePrime = 1;
	end	else if (num==16'd23593) begin
		AssumePrime = 1;
	end	else if (num==16'd23599) begin
		AssumePrime = 1;
	end	else if (num==16'd23603) begin
		AssumePrime = 1;
	end	else if (num==16'd23609) begin
		AssumePrime = 1;
	end	else if (num==16'd23623) begin
		AssumePrime = 1;
	end	else if (num==16'd23627) begin
		AssumePrime = 1;
	end	else if (num==16'd23629) begin
		AssumePrime = 1;
	end	else if (num==16'd23633) begin
		AssumePrime = 1;
	end	else if (num==16'd23663) begin
		AssumePrime = 1;
	end	else if (num==16'd23669) begin
		AssumePrime = 1;
	end	else if (num==16'd23671) begin
		AssumePrime = 1;
	end	else if (num==16'd23677) begin
		AssumePrime = 1;
	end	else if (num==16'd23687) begin
		AssumePrime = 1;
	end	else if (num==16'd23689) begin
		AssumePrime = 1;
	end	else if (num==16'd23719) begin
		AssumePrime = 1;
	end	else if (num==16'd23741) begin
		AssumePrime = 1;
	end	else if (num==16'd23743) begin
		AssumePrime = 1;
	end	else if (num==16'd23747) begin
		AssumePrime = 1;
	end	else if (num==16'd23753) begin
		AssumePrime = 1;
	end	else if (num==16'd23761) begin
		AssumePrime = 1;
	end	else if (num==16'd23767) begin
		AssumePrime = 1;
	end	else if (num==16'd23773) begin
		AssumePrime = 1;
	end	else if (num==16'd23789) begin
		AssumePrime = 1;
	end	else if (num==16'd23801) begin
		AssumePrime = 1;
	end	else if (num==16'd23813) begin
		AssumePrime = 1;
	end	else if (num==16'd23819) begin
		AssumePrime = 1;
	end	else if (num==16'd23827) begin
		AssumePrime = 1;
	end	else if (num==16'd23831) begin
		AssumePrime = 1;
	end	else if (num==16'd23833) begin
		AssumePrime = 1;
	end	else if (num==16'd23857) begin
		AssumePrime = 1;
	end	else if (num==16'd23869) begin
		AssumePrime = 1;
	end	else if (num==16'd23873) begin
		AssumePrime = 1;
	end	else if (num==16'd23879) begin
		AssumePrime = 1;
	end	else if (num==16'd23887) begin
		AssumePrime = 1;
	end	else if (num==16'd23893) begin
		AssumePrime = 1;
	end	else if (num==16'd23899) begin
		AssumePrime = 1;
	end	else if (num==16'd23909) begin
		AssumePrime = 1;
	end	else if (num==16'd23911) begin
		AssumePrime = 1;
	end	else if (num==16'd23917) begin
		AssumePrime = 1;
	end	else if (num==16'd23929) begin
		AssumePrime = 1;
	end	else if (num==16'd23957) begin
		AssumePrime = 1;
	end	else if (num==16'd23971) begin
		AssumePrime = 1;
	end	else if (num==16'd23977) begin
		AssumePrime = 1;
	end	else if (num==16'd23981) begin
		AssumePrime = 1;
	end	else if (num==16'd23993) begin
		AssumePrime = 1;
	end	else if (num==16'd24001) begin
		AssumePrime = 1;
	end	else if (num==16'd24007) begin
		AssumePrime = 1;
	end	else if (num==16'd24019) begin
		AssumePrime = 1;
	end	else if (num==16'd24023) begin
		AssumePrime = 1;
	end	else if (num==16'd24029) begin
		AssumePrime = 1;
	end	else if (num==16'd24043) begin
		AssumePrime = 1;
	end	else if (num==16'd24049) begin
		AssumePrime = 1;
	end	else if (num==16'd24061) begin
		AssumePrime = 1;
	end	else if (num==16'd24071) begin
		AssumePrime = 1;
	end	else if (num==16'd24077) begin
		AssumePrime = 1;
	end	else if (num==16'd24083) begin
		AssumePrime = 1;
	end	else if (num==16'd24091) begin
		AssumePrime = 1;
	end	else if (num==16'd24097) begin
		AssumePrime = 1;
	end	else if (num==16'd24103) begin
		AssumePrime = 1;
	end	else if (num==16'd24107) begin
		AssumePrime = 1;
	end	else if (num==16'd24109) begin
		AssumePrime = 1;
	end	else if (num==16'd24113) begin
		AssumePrime = 1;
	end	else if (num==16'd24121) begin
		AssumePrime = 1;
	end	else if (num==16'd24133) begin
		AssumePrime = 1;
	end	else if (num==16'd24137) begin
		AssumePrime = 1;
	end	else if (num==16'd24151) begin
		AssumePrime = 1;
	end	else if (num==16'd24169) begin
		AssumePrime = 1;
	end	else if (num==16'd24179) begin
		AssumePrime = 1;
	end	else if (num==16'd24181) begin
		AssumePrime = 1;
	end	else if (num==16'd24197) begin
		AssumePrime = 1;
	end	else if (num==16'd24203) begin
		AssumePrime = 1;
	end	else if (num==16'd24223) begin
		AssumePrime = 1;
	end	else if (num==16'd24229) begin
		AssumePrime = 1;
	end	else if (num==16'd24239) begin
		AssumePrime = 1;
	end	else if (num==16'd24247) begin
		AssumePrime = 1;
	end	else if (num==16'd24251) begin
		AssumePrime = 1;
	end	else if (num==16'd24281) begin
		AssumePrime = 1;
	end	else if (num==16'd24317) begin
		AssumePrime = 1;
	end	else if (num==16'd24329) begin
		AssumePrime = 1;
	end	else if (num==16'd24337) begin
		AssumePrime = 1;
	end	else if (num==16'd24359) begin
		AssumePrime = 1;
	end	else if (num==16'd24371) begin
		AssumePrime = 1;
	end	else if (num==16'd24373) begin
		AssumePrime = 1;
	end	else if (num==16'd24379) begin
		AssumePrime = 1;
	end	else if (num==16'd24391) begin
		AssumePrime = 1;
	end	else if (num==16'd24407) begin
		AssumePrime = 1;
	end	else if (num==16'd24413) begin
		AssumePrime = 1;
	end	else if (num==16'd24419) begin
		AssumePrime = 1;
	end	else if (num==16'd24421) begin
		AssumePrime = 1;
	end	else if (num==16'd24439) begin
		AssumePrime = 1;
	end	else if (num==16'd24443) begin
		AssumePrime = 1;
	end	else if (num==16'd24469) begin
		AssumePrime = 1;
	end	else if (num==16'd24473) begin
		AssumePrime = 1;
	end	else if (num==16'd24481) begin
		AssumePrime = 1;
	end	else if (num==16'd24499) begin
		AssumePrime = 1;
	end	else if (num==16'd24509) begin
		AssumePrime = 1;
	end	else if (num==16'd24517) begin
		AssumePrime = 1;
	end	else if (num==16'd24527) begin
		AssumePrime = 1;
	end	else if (num==16'd24533) begin
		AssumePrime = 1;
	end	else if (num==16'd24547) begin
		AssumePrime = 1;
	end	else if (num==16'd24551) begin
		AssumePrime = 1;
	end	else if (num==16'd24571) begin
		AssumePrime = 1;
	end	else if (num==16'd24593) begin
		AssumePrime = 1;
	end	else if (num==16'd24611) begin
		AssumePrime = 1;
	end	else if (num==16'd24623) begin
		AssumePrime = 1;
	end	else if (num==16'd24631) begin
		AssumePrime = 1;
	end	else if (num==16'd24659) begin
		AssumePrime = 1;
	end	else if (num==16'd24671) begin
		AssumePrime = 1;
	end	else if (num==16'd24677) begin
		AssumePrime = 1;
	end	else if (num==16'd24683) begin
		AssumePrime = 1;
	end	else if (num==16'd24691) begin
		AssumePrime = 1;
	end	else if (num==16'd24697) begin
		AssumePrime = 1;
	end	else if (num==16'd24709) begin
		AssumePrime = 1;
	end	else if (num==16'd24733) begin
		AssumePrime = 1;
	end	else if (num==16'd24749) begin
		AssumePrime = 1;
	end	else if (num==16'd24763) begin
		AssumePrime = 1;
	end	else if (num==16'd24767) begin
		AssumePrime = 1;
	end	else if (num==16'd24781) begin
		AssumePrime = 1;
	end	else if (num==16'd24793) begin
		AssumePrime = 1;
	end	else if (num==16'd24799) begin
		AssumePrime = 1;
	end	else if (num==16'd24809) begin
		AssumePrime = 1;
	end	else if (num==16'd24821) begin
		AssumePrime = 1;
	end	else if (num==16'd24841) begin
		AssumePrime = 1;
	end	else if (num==16'd24847) begin
		AssumePrime = 1;
	end	else if (num==16'd24851) begin
		AssumePrime = 1;
	end	else if (num==16'd24859) begin
		AssumePrime = 1;
	end	else if (num==16'd24877) begin
		AssumePrime = 1;
	end	else if (num==16'd24889) begin
		AssumePrime = 1;
	end	else if (num==16'd24907) begin
		AssumePrime = 1;
	end	else if (num==16'd24917) begin
		AssumePrime = 1;
	end	else if (num==16'd24919) begin
		AssumePrime = 1;
	end	else if (num==16'd24923) begin
		AssumePrime = 1;
	end	else if (num==16'd24943) begin
		AssumePrime = 1;
	end	else if (num==16'd24953) begin
		AssumePrime = 1;
	end	else if (num==16'd24967) begin
		AssumePrime = 1;
	end	else if (num==16'd24971) begin
		AssumePrime = 1;
	end	else if (num==16'd24977) begin
		AssumePrime = 1;
	end	else if (num==16'd24979) begin
		AssumePrime = 1;
	end	else if (num==16'd24989) begin
		AssumePrime = 1;
	end	else if (num==16'd25013) begin
		AssumePrime = 1;
	end	else if (num==16'd25031) begin
		AssumePrime = 1;
	end	else if (num==16'd25033) begin
		AssumePrime = 1;
	end	else if (num==16'd25037) begin
		AssumePrime = 1;
	end	else if (num==16'd25057) begin
		AssumePrime = 1;
	end	else if (num==16'd25073) begin
		AssumePrime = 1;
	end	else if (num==16'd25087) begin
		AssumePrime = 1;
	end	else if (num==16'd25097) begin
		AssumePrime = 1;
	end	else if (num==16'd25111) begin
		AssumePrime = 1;
	end	else if (num==16'd25117) begin
		AssumePrime = 1;
	end	else if (num==16'd25121) begin
		AssumePrime = 1;
	end	else if (num==16'd25127) begin
		AssumePrime = 1;
	end	else if (num==16'd25147) begin
		AssumePrime = 1;
	end	else if (num==16'd25153) begin
		AssumePrime = 1;
	end	else if (num==16'd25163) begin
		AssumePrime = 1;
	end	else if (num==16'd25169) begin
		AssumePrime = 1;
	end	else if (num==16'd25171) begin
		AssumePrime = 1;
	end	else if (num==16'd25183) begin
		AssumePrime = 1;
	end	else if (num==16'd25189) begin
		AssumePrime = 1;
	end	else if (num==16'd25219) begin
		AssumePrime = 1;
	end	else if (num==16'd25229) begin
		AssumePrime = 1;
	end	else if (num==16'd25237) begin
		AssumePrime = 1;
	end	else if (num==16'd25243) begin
		AssumePrime = 1;
	end	else if (num==16'd25247) begin
		AssumePrime = 1;
	end	else if (num==16'd25253) begin
		AssumePrime = 1;
	end	else if (num==16'd25261) begin
		AssumePrime = 1;
	end	else if (num==16'd25301) begin
		AssumePrime = 1;
	end	else if (num==16'd25303) begin
		AssumePrime = 1;
	end	else if (num==16'd25307) begin
		AssumePrime = 1;
	end	else if (num==16'd25309) begin
		AssumePrime = 1;
	end	else if (num==16'd25321) begin
		AssumePrime = 1;
	end	else if (num==16'd25339) begin
		AssumePrime = 1;
	end	else if (num==16'd25343) begin
		AssumePrime = 1;
	end	else if (num==16'd25349) begin
		AssumePrime = 1;
	end	else if (num==16'd25357) begin
		AssumePrime = 1;
	end	else if (num==16'd25367) begin
		AssumePrime = 1;
	end	else if (num==16'd25373) begin
		AssumePrime = 1;
	end	else if (num==16'd25391) begin
		AssumePrime = 1;
	end	else if (num==16'd25409) begin
		AssumePrime = 1;
	end	else if (num==16'd25411) begin
		AssumePrime = 1;
	end	else if (num==16'd25423) begin
		AssumePrime = 1;
	end	else if (num==16'd25439) begin
		AssumePrime = 1;
	end	else if (num==16'd25447) begin
		AssumePrime = 1;
	end	else if (num==16'd25453) begin
		AssumePrime = 1;
	end	else if (num==16'd25457) begin
		AssumePrime = 1;
	end	else if (num==16'd25463) begin
		AssumePrime = 1;
	end	else if (num==16'd25469) begin
		AssumePrime = 1;
	end	else if (num==16'd25471) begin
		AssumePrime = 1;
	end	else if (num==16'd25523) begin
		AssumePrime = 1;
	end	else if (num==16'd25537) begin
		AssumePrime = 1;
	end	else if (num==16'd25541) begin
		AssumePrime = 1;
	end	else if (num==16'd25561) begin
		AssumePrime = 1;
	end	else if (num==16'd25577) begin
		AssumePrime = 1;
	end	else if (num==16'd25579) begin
		AssumePrime = 1;
	end	else if (num==16'd25583) begin
		AssumePrime = 1;
	end	else if (num==16'd25589) begin
		AssumePrime = 1;
	end	else if (num==16'd25601) begin
		AssumePrime = 1;
	end	else if (num==16'd25603) begin
		AssumePrime = 1;
	end	else if (num==16'd25609) begin
		AssumePrime = 1;
	end	else if (num==16'd25621) begin
		AssumePrime = 1;
	end	else if (num==16'd25633) begin
		AssumePrime = 1;
	end	else if (num==16'd25639) begin
		AssumePrime = 1;
	end	else if (num==16'd25643) begin
		AssumePrime = 1;
	end	else if (num==16'd25657) begin
		AssumePrime = 1;
	end	else if (num==16'd25667) begin
		AssumePrime = 1;
	end	else if (num==16'd25673) begin
		AssumePrime = 1;
	end	else if (num==16'd25679) begin
		AssumePrime = 1;
	end	else if (num==16'd25693) begin
		AssumePrime = 1;
	end	else if (num==16'd25703) begin
		AssumePrime = 1;
	end	else if (num==16'd25717) begin
		AssumePrime = 1;
	end	else if (num==16'd25733) begin
		AssumePrime = 1;
	end	else if (num==16'd25741) begin
		AssumePrime = 1;
	end	else if (num==16'd25747) begin
		AssumePrime = 1;
	end	else if (num==16'd25759) begin
		AssumePrime = 1;
	end	else if (num==16'd25763) begin
		AssumePrime = 1;
	end	else if (num==16'd25771) begin
		AssumePrime = 1;
	end	else if (num==16'd25793) begin
		AssumePrime = 1;
	end	else if (num==16'd25799) begin
		AssumePrime = 1;
	end	else if (num==16'd25801) begin
		AssumePrime = 1;
	end	else if (num==16'd25819) begin
		AssumePrime = 1;
	end	else if (num==16'd25841) begin
		AssumePrime = 1;
	end	else if (num==16'd25847) begin
		AssumePrime = 1;
	end	else if (num==16'd25849) begin
		AssumePrime = 1;
	end	else if (num==16'd25867) begin
		AssumePrime = 1;
	end	else if (num==16'd25873) begin
		AssumePrime = 1;
	end	else if (num==16'd25889) begin
		AssumePrime = 1;
	end	else if (num==16'd25903) begin
		AssumePrime = 1;
	end	else if (num==16'd25913) begin
		AssumePrime = 1;
	end	else if (num==16'd25919) begin
		AssumePrime = 1;
	end	else if (num==16'd25931) begin
		AssumePrime = 1;
	end	else if (num==16'd25933) begin
		AssumePrime = 1;
	end	else if (num==16'd25939) begin
		AssumePrime = 1;
	end	else if (num==16'd25943) begin
		AssumePrime = 1;
	end	else if (num==16'd25951) begin
		AssumePrime = 1;
	end	else if (num==16'd25969) begin
		AssumePrime = 1;
	end	else if (num==16'd25981) begin
		AssumePrime = 1;
	end	else if (num==16'd25997) begin
		AssumePrime = 1;
	end	else if (num==16'd25999) begin
		AssumePrime = 1;
	end	else if (num==16'd26003) begin
		AssumePrime = 1;
	end	else if (num==16'd26017) begin
		AssumePrime = 1;
	end	else if (num==16'd26021) begin
		AssumePrime = 1;
	end	else if (num==16'd26029) begin
		AssumePrime = 1;
	end	else if (num==16'd26041) begin
		AssumePrime = 1;
	end	else if (num==16'd26053) begin
		AssumePrime = 1;
	end	else if (num==16'd26083) begin
		AssumePrime = 1;
	end	else if (num==16'd26099) begin
		AssumePrime = 1;
	end	else if (num==16'd26107) begin
		AssumePrime = 1;
	end	else if (num==16'd26111) begin
		AssumePrime = 1;
	end	else if (num==16'd26113) begin
		AssumePrime = 1;
	end	else if (num==16'd26119) begin
		AssumePrime = 1;
	end	else if (num==16'd26141) begin
		AssumePrime = 1;
	end	else if (num==16'd26153) begin
		AssumePrime = 1;
	end	else if (num==16'd26161) begin
		AssumePrime = 1;
	end	else if (num==16'd26171) begin
		AssumePrime = 1;
	end	else if (num==16'd26177) begin
		AssumePrime = 1;
	end	else if (num==16'd26183) begin
		AssumePrime = 1;
	end	else if (num==16'd26189) begin
		AssumePrime = 1;
	end	else if (num==16'd26203) begin
		AssumePrime = 1;
	end	else if (num==16'd26209) begin
		AssumePrime = 1;
	end	else if (num==16'd26227) begin
		AssumePrime = 1;
	end	else if (num==16'd26237) begin
		AssumePrime = 1;
	end	else if (num==16'd26249) begin
		AssumePrime = 1;
	end	else if (num==16'd26251) begin
		AssumePrime = 1;
	end	else if (num==16'd26261) begin
		AssumePrime = 1;
	end	else if (num==16'd26263) begin
		AssumePrime = 1;
	end	else if (num==16'd26267) begin
		AssumePrime = 1;
	end	else if (num==16'd26293) begin
		AssumePrime = 1;
	end	else if (num==16'd26297) begin
		AssumePrime = 1;
	end	else if (num==16'd26309) begin
		AssumePrime = 1;
	end	else if (num==16'd26317) begin
		AssumePrime = 1;
	end	else if (num==16'd26321) begin
		AssumePrime = 1;
	end	else if (num==16'd26339) begin
		AssumePrime = 1;
	end	else if (num==16'd26347) begin
		AssumePrime = 1;
	end	else if (num==16'd26357) begin
		AssumePrime = 1;
	end	else if (num==16'd26371) begin
		AssumePrime = 1;
	end	else if (num==16'd26387) begin
		AssumePrime = 1;
	end	else if (num==16'd26393) begin
		AssumePrime = 1;
	end	else if (num==16'd26399) begin
		AssumePrime = 1;
	end	else if (num==16'd26407) begin
		AssumePrime = 1;
	end	else if (num==16'd26417) begin
		AssumePrime = 1;
	end	else if (num==16'd26423) begin
		AssumePrime = 1;
	end	else if (num==16'd26431) begin
		AssumePrime = 1;
	end	else if (num==16'd26437) begin
		AssumePrime = 1;
	end	else if (num==16'd26449) begin
		AssumePrime = 1;
	end	else if (num==16'd26459) begin
		AssumePrime = 1;
	end	else if (num==16'd26479) begin
		AssumePrime = 1;
	end	else if (num==16'd26489) begin
		AssumePrime = 1;
	end	else if (num==16'd26497) begin
		AssumePrime = 1;
	end	else if (num==16'd26501) begin
		AssumePrime = 1;
	end	else if (num==16'd26513) begin
		AssumePrime = 1;
	end	else if (num==16'd26539) begin
		AssumePrime = 1;
	end	else if (num==16'd26557) begin
		AssumePrime = 1;
	end	else if (num==16'd26561) begin
		AssumePrime = 1;
	end	else if (num==16'd26573) begin
		AssumePrime = 1;
	end	else if (num==16'd26591) begin
		AssumePrime = 1;
	end	else if (num==16'd26597) begin
		AssumePrime = 1;
	end	else if (num==16'd26627) begin
		AssumePrime = 1;
	end	else if (num==16'd26633) begin
		AssumePrime = 1;
	end	else if (num==16'd26641) begin
		AssumePrime = 1;
	end	else if (num==16'd26647) begin
		AssumePrime = 1;
	end	else if (num==16'd26669) begin
		AssumePrime = 1;
	end	else if (num==16'd26681) begin
		AssumePrime = 1;
	end	else if (num==16'd26683) begin
		AssumePrime = 1;
	end	else if (num==16'd26687) begin
		AssumePrime = 1;
	end	else if (num==16'd26693) begin
		AssumePrime = 1;
	end	else if (num==16'd26699) begin
		AssumePrime = 1;
	end	else if (num==16'd26701) begin
		AssumePrime = 1;
	end	else if (num==16'd26711) begin
		AssumePrime = 1;
	end	else if (num==16'd26713) begin
		AssumePrime = 1;
	end	else if (num==16'd26717) begin
		AssumePrime = 1;
	end	else if (num==16'd26723) begin
		AssumePrime = 1;
	end	else if (num==16'd26729) begin
		AssumePrime = 1;
	end	else if (num==16'd26731) begin
		AssumePrime = 1;
	end	else if (num==16'd26737) begin
		AssumePrime = 1;
	end	else if (num==16'd26759) begin
		AssumePrime = 1;
	end	else if (num==16'd26777) begin
		AssumePrime = 1;
	end	else if (num==16'd26783) begin
		AssumePrime = 1;
	end	else if (num==16'd26801) begin
		AssumePrime = 1;
	end	else if (num==16'd26813) begin
		AssumePrime = 1;
	end	else if (num==16'd26821) begin
		AssumePrime = 1;
	end	else if (num==16'd26833) begin
		AssumePrime = 1;
	end	else if (num==16'd26839) begin
		AssumePrime = 1;
	end	else if (num==16'd26849) begin
		AssumePrime = 1;
	end	else if (num==16'd26861) begin
		AssumePrime = 1;
	end	else if (num==16'd26863) begin
		AssumePrime = 1;
	end	else if (num==16'd26879) begin
		AssumePrime = 1;
	end	else if (num==16'd26881) begin
		AssumePrime = 1;
	end	else if (num==16'd26891) begin
		AssumePrime = 1;
	end	else if (num==16'd26893) begin
		AssumePrime = 1;
	end	else if (num==16'd26903) begin
		AssumePrime = 1;
	end	else if (num==16'd26921) begin
		AssumePrime = 1;
	end	else if (num==16'd26927) begin
		AssumePrime = 1;
	end	else if (num==16'd26947) begin
		AssumePrime = 1;
	end	else if (num==16'd26951) begin
		AssumePrime = 1;
	end	else if (num==16'd26953) begin
		AssumePrime = 1;
	end	else if (num==16'd26959) begin
		AssumePrime = 1;
	end	else if (num==16'd26981) begin
		AssumePrime = 1;
	end	else if (num==16'd26987) begin
		AssumePrime = 1;
	end	else if (num==16'd26993) begin
		AssumePrime = 1;
	end	else if (num==16'd27011) begin
		AssumePrime = 1;
	end	else if (num==16'd27017) begin
		AssumePrime = 1;
	end	else if (num==16'd27031) begin
		AssumePrime = 1;
	end	else if (num==16'd27043) begin
		AssumePrime = 1;
	end	else if (num==16'd27059) begin
		AssumePrime = 1;
	end	else if (num==16'd27061) begin
		AssumePrime = 1;
	end	else if (num==16'd27067) begin
		AssumePrime = 1;
	end	else if (num==16'd27073) begin
		AssumePrime = 1;
	end	else if (num==16'd27077) begin
		AssumePrime = 1;
	end	else if (num==16'd27091) begin
		AssumePrime = 1;
	end	else if (num==16'd27103) begin
		AssumePrime = 1;
	end	else if (num==16'd27107) begin
		AssumePrime = 1;
	end	else if (num==16'd27109) begin
		AssumePrime = 1;
	end	else if (num==16'd27127) begin
		AssumePrime = 1;
	end	else if (num==16'd27143) begin
		AssumePrime = 1;
	end	else if (num==16'd27179) begin
		AssumePrime = 1;
	end	else if (num==16'd27191) begin
		AssumePrime = 1;
	end	else if (num==16'd27197) begin
		AssumePrime = 1;
	end	else if (num==16'd27211) begin
		AssumePrime = 1;
	end	else if (num==16'd27239) begin
		AssumePrime = 1;
	end	else if (num==16'd27241) begin
		AssumePrime = 1;
	end	else if (num==16'd27253) begin
		AssumePrime = 1;
	end	else if (num==16'd27259) begin
		AssumePrime = 1;
	end	else if (num==16'd27271) begin
		AssumePrime = 1;
	end	else if (num==16'd27277) begin
		AssumePrime = 1;
	end	else if (num==16'd27281) begin
		AssumePrime = 1;
	end	else if (num==16'd27283) begin
		AssumePrime = 1;
	end	else if (num==16'd27299) begin
		AssumePrime = 1;
	end	else if (num==16'd27329) begin
		AssumePrime = 1;
	end	else if (num==16'd27337) begin
		AssumePrime = 1;
	end	else if (num==16'd27361) begin
		AssumePrime = 1;
	end	else if (num==16'd27367) begin
		AssumePrime = 1;
	end	else if (num==16'd27397) begin
		AssumePrime = 1;
	end	else if (num==16'd27407) begin
		AssumePrime = 1;
	end	else if (num==16'd27409) begin
		AssumePrime = 1;
	end	else if (num==16'd27427) begin
		AssumePrime = 1;
	end	else if (num==16'd27431) begin
		AssumePrime = 1;
	end	else if (num==16'd27437) begin
		AssumePrime = 1;
	end	else if (num==16'd27449) begin
		AssumePrime = 1;
	end	else if (num==16'd27457) begin
		AssumePrime = 1;
	end	else if (num==16'd27479) begin
		AssumePrime = 1;
	end	else if (num==16'd27481) begin
		AssumePrime = 1;
	end	else if (num==16'd27487) begin
		AssumePrime = 1;
	end	else if (num==16'd27509) begin
		AssumePrime = 1;
	end	else if (num==16'd27527) begin
		AssumePrime = 1;
	end	else if (num==16'd27529) begin
		AssumePrime = 1;
	end	else if (num==16'd27539) begin
		AssumePrime = 1;
	end	else if (num==16'd27541) begin
		AssumePrime = 1;
	end	else if (num==16'd27551) begin
		AssumePrime = 1;
	end	else if (num==16'd27581) begin
		AssumePrime = 1;
	end	else if (num==16'd27583) begin
		AssumePrime = 1;
	end	else if (num==16'd27611) begin
		AssumePrime = 1;
	end	else if (num==16'd27617) begin
		AssumePrime = 1;
	end	else if (num==16'd27631) begin
		AssumePrime = 1;
	end	else if (num==16'd27647) begin
		AssumePrime = 1;
	end	else if (num==16'd27653) begin
		AssumePrime = 1;
	end	else if (num==16'd27673) begin
		AssumePrime = 1;
	end	else if (num==16'd27689) begin
		AssumePrime = 1;
	end	else if (num==16'd27691) begin
		AssumePrime = 1;
	end	else if (num==16'd27697) begin
		AssumePrime = 1;
	end	else if (num==16'd27701) begin
		AssumePrime = 1;
	end	else if (num==16'd27733) begin
		AssumePrime = 1;
	end	else if (num==16'd27737) begin
		AssumePrime = 1;
	end	else if (num==16'd27739) begin
		AssumePrime = 1;
	end	else if (num==16'd27743) begin
		AssumePrime = 1;
	end	else if (num==16'd27749) begin
		AssumePrime = 1;
	end	else if (num==16'd27751) begin
		AssumePrime = 1;
	end	else if (num==16'd27763) begin
		AssumePrime = 1;
	end	else if (num==16'd27767) begin
		AssumePrime = 1;
	end	else if (num==16'd27773) begin
		AssumePrime = 1;
	end	else if (num==16'd27779) begin
		AssumePrime = 1;
	end	else if (num==16'd27791) begin
		AssumePrime = 1;
	end	else if (num==16'd27793) begin
		AssumePrime = 1;
	end	else if (num==16'd27799) begin
		AssumePrime = 1;
	end	else if (num==16'd27803) begin
		AssumePrime = 1;
	end	else if (num==16'd27809) begin
		AssumePrime = 1;
	end	else if (num==16'd27817) begin
		AssumePrime = 1;
	end	else if (num==16'd27823) begin
		AssumePrime = 1;
	end	else if (num==16'd27827) begin
		AssumePrime = 1;
	end	else if (num==16'd27847) begin
		AssumePrime = 1;
	end	else if (num==16'd27851) begin
		AssumePrime = 1;
	end	else if (num==16'd27883) begin
		AssumePrime = 1;
	end	else if (num==16'd27893) begin
		AssumePrime = 1;
	end	else if (num==16'd27901) begin
		AssumePrime = 1;
	end	else if (num==16'd27917) begin
		AssumePrime = 1;
	end	else if (num==16'd27919) begin
		AssumePrime = 1;
	end	else if (num==16'd27941) begin
		AssumePrime = 1;
	end	else if (num==16'd27943) begin
		AssumePrime = 1;
	end	else if (num==16'd27947) begin
		AssumePrime = 1;
	end	else if (num==16'd27953) begin
		AssumePrime = 1;
	end	else if (num==16'd27961) begin
		AssumePrime = 1;
	end	else if (num==16'd27967) begin
		AssumePrime = 1;
	end	else if (num==16'd27983) begin
		AssumePrime = 1;
	end	else if (num==16'd27997) begin
		AssumePrime = 1;
	end	else if (num==16'd28001) begin
		AssumePrime = 1;
	end	else if (num==16'd28019) begin
		AssumePrime = 1;
	end	else if (num==16'd28027) begin
		AssumePrime = 1;
	end	else if (num==16'd28031) begin
		AssumePrime = 1;
	end	else if (num==16'd28051) begin
		AssumePrime = 1;
	end	else if (num==16'd28057) begin
		AssumePrime = 1;
	end	else if (num==16'd28069) begin
		AssumePrime = 1;
	end	else if (num==16'd28081) begin
		AssumePrime = 1;
	end	else if (num==16'd28087) begin
		AssumePrime = 1;
	end	else if (num==16'd28097) begin
		AssumePrime = 1;
	end	else if (num==16'd28099) begin
		AssumePrime = 1;
	end	else if (num==16'd28109) begin
		AssumePrime = 1;
	end	else if (num==16'd28111) begin
		AssumePrime = 1;
	end	else if (num==16'd28123) begin
		AssumePrime = 1;
	end	else if (num==16'd28151) begin
		AssumePrime = 1;
	end	else if (num==16'd28163) begin
		AssumePrime = 1;
	end	else if (num==16'd28181) begin
		AssumePrime = 1;
	end	else if (num==16'd28183) begin
		AssumePrime = 1;
	end	else if (num==16'd28201) begin
		AssumePrime = 1;
	end	else if (num==16'd28211) begin
		AssumePrime = 1;
	end	else if (num==16'd28219) begin
		AssumePrime = 1;
	end	else if (num==16'd28229) begin
		AssumePrime = 1;
	end	else if (num==16'd28277) begin
		AssumePrime = 1;
	end	else if (num==16'd28279) begin
		AssumePrime = 1;
	end	else if (num==16'd28283) begin
		AssumePrime = 1;
	end	else if (num==16'd28289) begin
		AssumePrime = 1;
	end	else if (num==16'd28297) begin
		AssumePrime = 1;
	end	else if (num==16'd28307) begin
		AssumePrime = 1;
	end	else if (num==16'd28309) begin
		AssumePrime = 1;
	end	else if (num==16'd28319) begin
		AssumePrime = 1;
	end	else if (num==16'd28349) begin
		AssumePrime = 1;
	end	else if (num==16'd28351) begin
		AssumePrime = 1;
	end	else if (num==16'd28387) begin
		AssumePrime = 1;
	end	else if (num==16'd28393) begin
		AssumePrime = 1;
	end	else if (num==16'd28403) begin
		AssumePrime = 1;
	end	else if (num==16'd28409) begin
		AssumePrime = 1;
	end	else if (num==16'd28411) begin
		AssumePrime = 1;
	end	else if (num==16'd28429) begin
		AssumePrime = 1;
	end	else if (num==16'd28433) begin
		AssumePrime = 1;
	end	else if (num==16'd28439) begin
		AssumePrime = 1;
	end	else if (num==16'd28447) begin
		AssumePrime = 1;
	end	else if (num==16'd28463) begin
		AssumePrime = 1;
	end	else if (num==16'd28477) begin
		AssumePrime = 1;
	end	else if (num==16'd28493) begin
		AssumePrime = 1;
	end	else if (num==16'd28499) begin
		AssumePrime = 1;
	end	else if (num==16'd28513) begin
		AssumePrime = 1;
	end	else if (num==16'd28517) begin
		AssumePrime = 1;
	end	else if (num==16'd28537) begin
		AssumePrime = 1;
	end	else if (num==16'd28541) begin
		AssumePrime = 1;
	end	else if (num==16'd28547) begin
		AssumePrime = 1;
	end	else if (num==16'd28549) begin
		AssumePrime = 1;
	end	else if (num==16'd28559) begin
		AssumePrime = 1;
	end	else if (num==16'd28571) begin
		AssumePrime = 1;
	end	else if (num==16'd28573) begin
		AssumePrime = 1;
	end	else if (num==16'd28579) begin
		AssumePrime = 1;
	end	else if (num==16'd28591) begin
		AssumePrime = 1;
	end	else if (num==16'd28597) begin
		AssumePrime = 1;
	end	else if (num==16'd28603) begin
		AssumePrime = 1;
	end	else if (num==16'd28607) begin
		AssumePrime = 1;
	end	else if (num==16'd28619) begin
		AssumePrime = 1;
	end	else if (num==16'd28621) begin
		AssumePrime = 1;
	end	else if (num==16'd28627) begin
		AssumePrime = 1;
	end	else if (num==16'd28631) begin
		AssumePrime = 1;
	end	else if (num==16'd28643) begin
		AssumePrime = 1;
	end	else if (num==16'd28649) begin
		AssumePrime = 1;
	end	else if (num==16'd28657) begin
		AssumePrime = 1;
	end	else if (num==16'd28661) begin
		AssumePrime = 1;
	end	else if (num==16'd28663) begin
		AssumePrime = 1;
	end	else if (num==16'd28669) begin
		AssumePrime = 1;
	end	else if (num==16'd28687) begin
		AssumePrime = 1;
	end	else if (num==16'd28697) begin
		AssumePrime = 1;
	end	else if (num==16'd28703) begin
		AssumePrime = 1;
	end	else if (num==16'd28711) begin
		AssumePrime = 1;
	end	else if (num==16'd28723) begin
		AssumePrime = 1;
	end	else if (num==16'd28729) begin
		AssumePrime = 1;
	end	else if (num==16'd28751) begin
		AssumePrime = 1;
	end	else if (num==16'd28753) begin
		AssumePrime = 1;
	end	else if (num==16'd28759) begin
		AssumePrime = 1;
	end	else if (num==16'd28771) begin
		AssumePrime = 1;
	end	else if (num==16'd28789) begin
		AssumePrime = 1;
	end	else if (num==16'd28793) begin
		AssumePrime = 1;
	end	else if (num==16'd28807) begin
		AssumePrime = 1;
	end	else if (num==16'd28813) begin
		AssumePrime = 1;
	end	else if (num==16'd28817) begin
		AssumePrime = 1;
	end	else if (num==16'd28837) begin
		AssumePrime = 1;
	end	else if (num==16'd28843) begin
		AssumePrime = 1;
	end	else if (num==16'd28859) begin
		AssumePrime = 1;
	end	else if (num==16'd28867) begin
		AssumePrime = 1;
	end	else if (num==16'd28871) begin
		AssumePrime = 1;
	end	else if (num==16'd28879) begin
		AssumePrime = 1;
	end	else if (num==16'd28901) begin
		AssumePrime = 1;
	end	else if (num==16'd28909) begin
		AssumePrime = 1;
	end	else if (num==16'd28921) begin
		AssumePrime = 1;
	end	else if (num==16'd28927) begin
		AssumePrime = 1;
	end	else if (num==16'd28933) begin
		AssumePrime = 1;
	end	else if (num==16'd28949) begin
		AssumePrime = 1;
	end	else if (num==16'd28961) begin
		AssumePrime = 1;
	end	else if (num==16'd28979) begin
		AssumePrime = 1;
	end	else if (num==16'd29009) begin
		AssumePrime = 1;
	end	else if (num==16'd29017) begin
		AssumePrime = 1;
	end	else if (num==16'd29021) begin
		AssumePrime = 1;
	end	else if (num==16'd29023) begin
		AssumePrime = 1;
	end	else if (num==16'd29027) begin
		AssumePrime = 1;
	end	else if (num==16'd29033) begin
		AssumePrime = 1;
	end	else if (num==16'd29059) begin
		AssumePrime = 1;
	end	else if (num==16'd29063) begin
		AssumePrime = 1;
	end	else if (num==16'd29077) begin
		AssumePrime = 1;
	end	else if (num==16'd29101) begin
		AssumePrime = 1;
	end	else if (num==16'd29123) begin
		AssumePrime = 1;
	end	else if (num==16'd29129) begin
		AssumePrime = 1;
	end	else if (num==16'd29131) begin
		AssumePrime = 1;
	end	else if (num==16'd29137) begin
		AssumePrime = 1;
	end	else if (num==16'd29147) begin
		AssumePrime = 1;
	end	else if (num==16'd29153) begin
		AssumePrime = 1;
	end	else if (num==16'd29167) begin
		AssumePrime = 1;
	end	else if (num==16'd29173) begin
		AssumePrime = 1;
	end	else if (num==16'd29179) begin
		AssumePrime = 1;
	end	else if (num==16'd29191) begin
		AssumePrime = 1;
	end	else if (num==16'd29201) begin
		AssumePrime = 1;
	end	else if (num==16'd29207) begin
		AssumePrime = 1;
	end	else if (num==16'd29209) begin
		AssumePrime = 1;
	end	else if (num==16'd29221) begin
		AssumePrime = 1;
	end	else if (num==16'd29231) begin
		AssumePrime = 1;
	end	else if (num==16'd29243) begin
		AssumePrime = 1;
	end	else if (num==16'd29251) begin
		AssumePrime = 1;
	end	else if (num==16'd29269) begin
		AssumePrime = 1;
	end	else if (num==16'd29287) begin
		AssumePrime = 1;
	end	else if (num==16'd29297) begin
		AssumePrime = 1;
	end	else if (num==16'd29303) begin
		AssumePrime = 1;
	end	else if (num==16'd29311) begin
		AssumePrime = 1;
	end	else if (num==16'd29327) begin
		AssumePrime = 1;
	end	else if (num==16'd29333) begin
		AssumePrime = 1;
	end	else if (num==16'd29339) begin
		AssumePrime = 1;
	end	else if (num==16'd29347) begin
		AssumePrime = 1;
	end	else if (num==16'd29363) begin
		AssumePrime = 1;
	end	else if (num==16'd29383) begin
		AssumePrime = 1;
	end	else if (num==16'd29387) begin
		AssumePrime = 1;
	end	else if (num==16'd29389) begin
		AssumePrime = 1;
	end	else if (num==16'd29399) begin
		AssumePrime = 1;
	end	else if (num==16'd29401) begin
		AssumePrime = 1;
	end	else if (num==16'd29411) begin
		AssumePrime = 1;
	end	else if (num==16'd29423) begin
		AssumePrime = 1;
	end	else if (num==16'd29429) begin
		AssumePrime = 1;
	end	else if (num==16'd29437) begin
		AssumePrime = 1;
	end	else if (num==16'd29443) begin
		AssumePrime = 1;
	end	else if (num==16'd29453) begin
		AssumePrime = 1;
	end	else if (num==16'd29473) begin
		AssumePrime = 1;
	end	else if (num==16'd29483) begin
		AssumePrime = 1;
	end	else if (num==16'd29501) begin
		AssumePrime = 1;
	end	else if (num==16'd29527) begin
		AssumePrime = 1;
	end	else if (num==16'd29531) begin
		AssumePrime = 1;
	end	else if (num==16'd29537) begin
		AssumePrime = 1;
	end	else if (num==16'd29567) begin
		AssumePrime = 1;
	end	else if (num==16'd29569) begin
		AssumePrime = 1;
	end	else if (num==16'd29573) begin
		AssumePrime = 1;
	end	else if (num==16'd29581) begin
		AssumePrime = 1;
	end	else if (num==16'd29587) begin
		AssumePrime = 1;
	end	else if (num==16'd29599) begin
		AssumePrime = 1;
	end	else if (num==16'd29611) begin
		AssumePrime = 1;
	end	else if (num==16'd29629) begin
		AssumePrime = 1;
	end	else if (num==16'd29633) begin
		AssumePrime = 1;
	end	else if (num==16'd29641) begin
		AssumePrime = 1;
	end	else if (num==16'd29663) begin
		AssumePrime = 1;
	end	else if (num==16'd29669) begin
		AssumePrime = 1;
	end	else if (num==16'd29671) begin
		AssumePrime = 1;
	end	else if (num==16'd29683) begin
		AssumePrime = 1;
	end	else if (num==16'd29717) begin
		AssumePrime = 1;
	end	else if (num==16'd29723) begin
		AssumePrime = 1;
	end	else if (num==16'd29741) begin
		AssumePrime = 1;
	end	else if (num==16'd29753) begin
		AssumePrime = 1;
	end	else if (num==16'd29759) begin
		AssumePrime = 1;
	end	else if (num==16'd29761) begin
		AssumePrime = 1;
	end	else if (num==16'd29789) begin
		AssumePrime = 1;
	end	else if (num==16'd29803) begin
		AssumePrime = 1;
	end	else if (num==16'd29819) begin
		AssumePrime = 1;
	end	else if (num==16'd29833) begin
		AssumePrime = 1;
	end	else if (num==16'd29837) begin
		AssumePrime = 1;
	end	else if (num==16'd29851) begin
		AssumePrime = 1;
	end	else if (num==16'd29863) begin
		AssumePrime = 1;
	end	else if (num==16'd29867) begin
		AssumePrime = 1;
	end	else if (num==16'd29873) begin
		AssumePrime = 1;
	end	else if (num==16'd29879) begin
		AssumePrime = 1;
	end	else if (num==16'd29881) begin
		AssumePrime = 1;
	end	else if (num==16'd29917) begin
		AssumePrime = 1;
	end	else if (num==16'd29921) begin
		AssumePrime = 1;
	end	else if (num==16'd29927) begin
		AssumePrime = 1;
	end	else if (num==16'd29947) begin
		AssumePrime = 1;
	end	else if (num==16'd29959) begin
		AssumePrime = 1;
	end	else if (num==16'd29983) begin
		AssumePrime = 1;
	end	else if (num==16'd29989) begin
		AssumePrime = 1;
	end	else if (num==16'd30011) begin
		AssumePrime = 1;
	end	else if (num==16'd30013) begin
		AssumePrime = 1;
	end	else if (num==16'd30029) begin
		AssumePrime = 1;
	end	else if (num==16'd30047) begin
		AssumePrime = 1;
	end	else if (num==16'd30059) begin
		AssumePrime = 1;
	end	else if (num==16'd30071) begin
		AssumePrime = 1;
	end	else if (num==16'd30089) begin
		AssumePrime = 1;
	end	else if (num==16'd30091) begin
		AssumePrime = 1;
	end	else if (num==16'd30097) begin
		AssumePrime = 1;
	end	else if (num==16'd30103) begin
		AssumePrime = 1;
	end	else if (num==16'd30109) begin
		AssumePrime = 1;
	end	else if (num==16'd30113) begin
		AssumePrime = 1;
	end	else if (num==16'd30119) begin
		AssumePrime = 1;
	end	else if (num==16'd30133) begin
		AssumePrime = 1;
	end	else if (num==16'd30137) begin
		AssumePrime = 1;
	end	else if (num==16'd30139) begin
		AssumePrime = 1;
	end	else if (num==16'd30161) begin
		AssumePrime = 1;
	end	else if (num==16'd30169) begin
		AssumePrime = 1;
	end	else if (num==16'd30181) begin
		AssumePrime = 1;
	end	else if (num==16'd30187) begin
		AssumePrime = 1;
	end	else if (num==16'd30197) begin
		AssumePrime = 1;
	end	else if (num==16'd30203) begin
		AssumePrime = 1;
	end	else if (num==16'd30211) begin
		AssumePrime = 1;
	end	else if (num==16'd30223) begin
		AssumePrime = 1;
	end	else if (num==16'd30241) begin
		AssumePrime = 1;
	end	else if (num==16'd30253) begin
		AssumePrime = 1;
	end	else if (num==16'd30259) begin
		AssumePrime = 1;
	end	else if (num==16'd30269) begin
		AssumePrime = 1;
	end	else if (num==16'd30271) begin
		AssumePrime = 1;
	end	else if (num==16'd30293) begin
		AssumePrime = 1;
	end	else if (num==16'd30307) begin
		AssumePrime = 1;
	end	else if (num==16'd30313) begin
		AssumePrime = 1;
	end	else if (num==16'd30319) begin
		AssumePrime = 1;
	end	else if (num==16'd30323) begin
		AssumePrime = 1;
	end	else if (num==16'd30341) begin
		AssumePrime = 1;
	end	else if (num==16'd30347) begin
		AssumePrime = 1;
	end	else if (num==16'd30367) begin
		AssumePrime = 1;
	end	else if (num==16'd30389) begin
		AssumePrime = 1;
	end	else if (num==16'd30391) begin
		AssumePrime = 1;
	end	else if (num==16'd30403) begin
		AssumePrime = 1;
	end	else if (num==16'd30427) begin
		AssumePrime = 1;
	end	else if (num==16'd30431) begin
		AssumePrime = 1;
	end	else if (num==16'd30449) begin
		AssumePrime = 1;
	end	else if (num==16'd30467) begin
		AssumePrime = 1;
	end	else if (num==16'd30469) begin
		AssumePrime = 1;
	end	else if (num==16'd30491) begin
		AssumePrime = 1;
	end	else if (num==16'd30493) begin
		AssumePrime = 1;
	end	else if (num==16'd30497) begin
		AssumePrime = 1;
	end	else if (num==16'd30509) begin
		AssumePrime = 1;
	end	else if (num==16'd30517) begin
		AssumePrime = 1;
	end	else if (num==16'd30529) begin
		AssumePrime = 1;
	end	else if (num==16'd30539) begin
		AssumePrime = 1;
	end	else if (num==16'd30553) begin
		AssumePrime = 1;
	end	else if (num==16'd30557) begin
		AssumePrime = 1;
	end	else if (num==16'd30559) begin
		AssumePrime = 1;
	end	else if (num==16'd30577) begin
		AssumePrime = 1;
	end	else if (num==16'd30593) begin
		AssumePrime = 1;
	end	else if (num==16'd30631) begin
		AssumePrime = 1;
	end	else if (num==16'd30637) begin
		AssumePrime = 1;
	end	else if (num==16'd30643) begin
		AssumePrime = 1;
	end	else if (num==16'd30649) begin
		AssumePrime = 1;
	end	else if (num==16'd30661) begin
		AssumePrime = 1;
	end	else if (num==16'd30671) begin
		AssumePrime = 1;
	end	else if (num==16'd30677) begin
		AssumePrime = 1;
	end	else if (num==16'd30689) begin
		AssumePrime = 1;
	end	else if (num==16'd30697) begin
		AssumePrime = 1;
	end	else if (num==16'd30703) begin
		AssumePrime = 1;
	end	else if (num==16'd30707) begin
		AssumePrime = 1;
	end	else if (num==16'd30713) begin
		AssumePrime = 1;
	end	else if (num==16'd30727) begin
		AssumePrime = 1;
	end	else if (num==16'd30757) begin
		AssumePrime = 1;
	end	else if (num==16'd30763) begin
		AssumePrime = 1;
	end	else if (num==16'd30773) begin
		AssumePrime = 1;
	end	else if (num==16'd30781) begin
		AssumePrime = 1;
	end	else if (num==16'd30803) begin
		AssumePrime = 1;
	end	else if (num==16'd30809) begin
		AssumePrime = 1;
	end	else if (num==16'd30817) begin
		AssumePrime = 1;
	end	else if (num==16'd30829) begin
		AssumePrime = 1;
	end	else if (num==16'd30839) begin
		AssumePrime = 1;
	end	else if (num==16'd30841) begin
		AssumePrime = 1;
	end	else if (num==16'd30851) begin
		AssumePrime = 1;
	end	else if (num==16'd30853) begin
		AssumePrime = 1;
	end	else if (num==16'd30859) begin
		AssumePrime = 1;
	end	else if (num==16'd30869) begin
		AssumePrime = 1;
	end	else if (num==16'd30871) begin
		AssumePrime = 1;
	end	else if (num==16'd30881) begin
		AssumePrime = 1;
	end	else if (num==16'd30893) begin
		AssumePrime = 1;
	end	else if (num==16'd30911) begin
		AssumePrime = 1;
	end	else if (num==16'd30931) begin
		AssumePrime = 1;
	end	else if (num==16'd30937) begin
		AssumePrime = 1;
	end	else if (num==16'd30941) begin
		AssumePrime = 1;
	end	else if (num==16'd30949) begin
		AssumePrime = 1;
	end	else if (num==16'd30971) begin
		AssumePrime = 1;
	end	else if (num==16'd30977) begin
		AssumePrime = 1;
	end	else if (num==16'd30983) begin
		AssumePrime = 1;
	end	else if (num==16'd31013) begin
		AssumePrime = 1;
	end	else if (num==16'd31019) begin
		AssumePrime = 1;
	end	else if (num==16'd31033) begin
		AssumePrime = 1;
	end	else if (num==16'd31039) begin
		AssumePrime = 1;
	end	else if (num==16'd31051) begin
		AssumePrime = 1;
	end	else if (num==16'd31063) begin
		AssumePrime = 1;
	end	else if (num==16'd31069) begin
		AssumePrime = 1;
	end	else if (num==16'd31079) begin
		AssumePrime = 1;
	end	else if (num==16'd31081) begin
		AssumePrime = 1;
	end	else if (num==16'd31091) begin
		AssumePrime = 1;
	end	else if (num==16'd31121) begin
		AssumePrime = 1;
	end	else if (num==16'd31123) begin
		AssumePrime = 1;
	end	else if (num==16'd31139) begin
		AssumePrime = 1;
	end	else if (num==16'd31147) begin
		AssumePrime = 1;
	end	else if (num==16'd31151) begin
		AssumePrime = 1;
	end	else if (num==16'd31153) begin
		AssumePrime = 1;
	end	else if (num==16'd31159) begin
		AssumePrime = 1;
	end	else if (num==16'd31177) begin
		AssumePrime = 1;
	end	else if (num==16'd31181) begin
		AssumePrime = 1;
	end	else if (num==16'd31183) begin
		AssumePrime = 1;
	end	else if (num==16'd31189) begin
		AssumePrime = 1;
	end	else if (num==16'd31193) begin
		AssumePrime = 1;
	end	else if (num==16'd31219) begin
		AssumePrime = 1;
	end	else if (num==16'd31223) begin
		AssumePrime = 1;
	end	else if (num==16'd31231) begin
		AssumePrime = 1;
	end	else if (num==16'd31237) begin
		AssumePrime = 1;
	end	else if (num==16'd31247) begin
		AssumePrime = 1;
	end	else if (num==16'd31249) begin
		AssumePrime = 1;
	end	else if (num==16'd31253) begin
		AssumePrime = 1;
	end	else if (num==16'd31259) begin
		AssumePrime = 1;
	end	else if (num==16'd31267) begin
		AssumePrime = 1;
	end	else if (num==16'd31271) begin
		AssumePrime = 1;
	end	else if (num==16'd31277) begin
		AssumePrime = 1;
	end	else if (num==16'd31307) begin
		AssumePrime = 1;
	end	else if (num==16'd31319) begin
		AssumePrime = 1;
	end	else if (num==16'd31321) begin
		AssumePrime = 1;
	end	else if (num==16'd31327) begin
		AssumePrime = 1;
	end	else if (num==16'd31333) begin
		AssumePrime = 1;
	end	else if (num==16'd31337) begin
		AssumePrime = 1;
	end	else if (num==16'd31357) begin
		AssumePrime = 1;
	end	else if (num==16'd31379) begin
		AssumePrime = 1;
	end	else if (num==16'd31387) begin
		AssumePrime = 1;
	end	else if (num==16'd31391) begin
		AssumePrime = 1;
	end	else if (num==16'd31393) begin
		AssumePrime = 1;
	end	else if (num==16'd31397) begin
		AssumePrime = 1;
	end	else if (num==16'd31469) begin
		AssumePrime = 1;
	end	else if (num==16'd31477) begin
		AssumePrime = 1;
	end	else if (num==16'd31481) begin
		AssumePrime = 1;
	end	else if (num==16'd31489) begin
		AssumePrime = 1;
	end	else if (num==16'd31511) begin
		AssumePrime = 1;
	end	else if (num==16'd31513) begin
		AssumePrime = 1;
	end	else if (num==16'd31517) begin
		AssumePrime = 1;
	end	else if (num==16'd31531) begin
		AssumePrime = 1;
	end	else if (num==16'd31541) begin
		AssumePrime = 1;
	end	else if (num==16'd31543) begin
		AssumePrime = 1;
	end	else if (num==16'd31547) begin
		AssumePrime = 1;
	end	else if (num==16'd31567) begin
		AssumePrime = 1;
	end	else if (num==16'd31573) begin
		AssumePrime = 1;
	end	else if (num==16'd31583) begin
		AssumePrime = 1;
	end	else if (num==16'd31601) begin
		AssumePrime = 1;
	end	else if (num==16'd31607) begin
		AssumePrime = 1;
	end	else if (num==16'd31627) begin
		AssumePrime = 1;
	end	else if (num==16'd31643) begin
		AssumePrime = 1;
	end	else if (num==16'd31649) begin
		AssumePrime = 1;
	end	else if (num==16'd31657) begin
		AssumePrime = 1;
	end	else if (num==16'd31663) begin
		AssumePrime = 1;
	end	else if (num==16'd31667) begin
		AssumePrime = 1;
	end	else if (num==16'd31687) begin
		AssumePrime = 1;
	end	else if (num==16'd31699) begin
		AssumePrime = 1;
	end	else if (num==16'd31721) begin
		AssumePrime = 1;
	end	else if (num==16'd31723) begin
		AssumePrime = 1;
	end	else if (num==16'd31727) begin
		AssumePrime = 1;
	end	else if (num==16'd31729) begin
		AssumePrime = 1;
	end	else if (num==16'd31741) begin
		AssumePrime = 1;
	end	else if (num==16'd31751) begin
		AssumePrime = 1;
	end	else if (num==16'd31769) begin
		AssumePrime = 1;
	end	else if (num==16'd31771) begin
		AssumePrime = 1;
	end	else if (num==16'd31793) begin
		AssumePrime = 1;
	end	else if (num==16'd31799) begin
		AssumePrime = 1;
	end	else if (num==16'd31817) begin
		AssumePrime = 1;
	end	else if (num==16'd31847) begin
		AssumePrime = 1;
	end	else if (num==16'd31849) begin
		AssumePrime = 1;
	end	else if (num==16'd31859) begin
		AssumePrime = 1;
	end	else if (num==16'd31873) begin
		AssumePrime = 1;
	end	else if (num==16'd31883) begin
		AssumePrime = 1;
	end	else if (num==16'd31891) begin
		AssumePrime = 1;
	end	else if (num==16'd31907) begin
		AssumePrime = 1;
	end	else if (num==16'd31957) begin
		AssumePrime = 1;
	end	else if (num==16'd31963) begin
		AssumePrime = 1;
	end	else if (num==16'd31973) begin
		AssumePrime = 1;
	end	else if (num==16'd31981) begin
		AssumePrime = 1;
	end	else if (num==16'd31991) begin
		AssumePrime = 1;
	end	else if (num==16'd32003) begin
		AssumePrime = 1;
	end	else if (num==16'd32009) begin
		AssumePrime = 1;
	end	else if (num==16'd32027) begin
		AssumePrime = 1;
	end	else if (num==16'd32029) begin
		AssumePrime = 1;
	end	else if (num==16'd32051) begin
		AssumePrime = 1;
	end	else if (num==16'd32057) begin
		AssumePrime = 1;
	end	else if (num==16'd32059) begin
		AssumePrime = 1;
	end	else if (num==16'd32063) begin
		AssumePrime = 1;
	end	else if (num==16'd32069) begin
		AssumePrime = 1;
	end	else if (num==16'd32077) begin
		AssumePrime = 1;
	end	else if (num==16'd32083) begin
		AssumePrime = 1;
	end	else if (num==16'd32089) begin
		AssumePrime = 1;
	end	else if (num==16'd32099) begin
		AssumePrime = 1;
	end	else if (num==16'd32117) begin
		AssumePrime = 1;
	end	else if (num==16'd32119) begin
		AssumePrime = 1;
	end	else if (num==16'd32141) begin
		AssumePrime = 1;
	end	else if (num==16'd32143) begin
		AssumePrime = 1;
	end	else if (num==16'd32159) begin
		AssumePrime = 1;
	end	else if (num==16'd32173) begin
		AssumePrime = 1;
	end	else if (num==16'd32183) begin
		AssumePrime = 1;
	end	else if (num==16'd32189) begin
		AssumePrime = 1;
	end	else if (num==16'd32191) begin
		AssumePrime = 1;
	end	else if (num==16'd32203) begin
		AssumePrime = 1;
	end	else if (num==16'd32213) begin
		AssumePrime = 1;
	end	else if (num==16'd32233) begin
		AssumePrime = 1;
	end	else if (num==16'd32237) begin
		AssumePrime = 1;
	end	else if (num==16'd32251) begin
		AssumePrime = 1;
	end	else if (num==16'd32257) begin
		AssumePrime = 1;
	end	else if (num==16'd32261) begin
		AssumePrime = 1;
	end	else if (num==16'd32297) begin
		AssumePrime = 1;
	end	else if (num==16'd32299) begin
		AssumePrime = 1;
	end	else if (num==16'd32303) begin
		AssumePrime = 1;
	end	else if (num==16'd32309) begin
		AssumePrime = 1;
	end	else if (num==16'd32321) begin
		AssumePrime = 1;
	end	else if (num==16'd32323) begin
		AssumePrime = 1;
	end	else if (num==16'd32327) begin
		AssumePrime = 1;
	end	else if (num==16'd32341) begin
		AssumePrime = 1;
	end	else if (num==16'd32353) begin
		AssumePrime = 1;
	end	else if (num==16'd32359) begin
		AssumePrime = 1;
	end	else if (num==16'd32363) begin
		AssumePrime = 1;
	end	else if (num==16'd32369) begin
		AssumePrime = 1;
	end	else if (num==16'd32371) begin
		AssumePrime = 1;
	end	else if (num==16'd32377) begin
		AssumePrime = 1;
	end	else if (num==16'd32381) begin
		AssumePrime = 1;
	end	else if (num==16'd32401) begin
		AssumePrime = 1;
	end	else if (num==16'd32411) begin
		AssumePrime = 1;
	end	else if (num==16'd32413) begin
		AssumePrime = 1;
	end	else if (num==16'd32423) begin
		AssumePrime = 1;
	end	else if (num==16'd32429) begin
		AssumePrime = 1;
	end	else if (num==16'd32441) begin
		AssumePrime = 1;
	end	else if (num==16'd32443) begin
		AssumePrime = 1;
	end	else if (num==16'd32467) begin
		AssumePrime = 1;
	end	else if (num==16'd32479) begin
		AssumePrime = 1;
	end	else if (num==16'd32491) begin
		AssumePrime = 1;
	end	else if (num==16'd32497) begin
		AssumePrime = 1;
	end	else if (num==16'd32503) begin
		AssumePrime = 1;
	end	else if (num==16'd32507) begin
		AssumePrime = 1;
	end	else if (num==16'd32531) begin
		AssumePrime = 1;
	end	else if (num==16'd32533) begin
		AssumePrime = 1;
	end	else if (num==16'd32537) begin
		AssumePrime = 1;
	end	else if (num==16'd32561) begin
		AssumePrime = 1;
	end	else if (num==16'd32563) begin
		AssumePrime = 1;
	end	else if (num==16'd32569) begin
		AssumePrime = 1;
	end	else if (num==16'd32573) begin
		AssumePrime = 1;
	end	else if (num==16'd32579) begin
		AssumePrime = 1;
	end	else if (num==16'd32587) begin
		AssumePrime = 1;
	end	else if (num==16'd32603) begin
		AssumePrime = 1;
	end	else if (num==16'd32609) begin
		AssumePrime = 1;
	end	else if (num==16'd32611) begin
		AssumePrime = 1;
	end	else if (num==16'd32621) begin
		AssumePrime = 1;
	end	else if (num==16'd32633) begin
		AssumePrime = 1;
	end	else if (num==16'd32647) begin
		AssumePrime = 1;
	end	else if (num==16'd32653) begin
		AssumePrime = 1;
	end	else if (num==16'd32687) begin
		AssumePrime = 1;
	end	else if (num==16'd32693) begin
		AssumePrime = 1;
	end	else if (num==16'd32707) begin
		AssumePrime = 1;
	end	else if (num==16'd32713) begin
		AssumePrime = 1;
	end	else if (num==16'd32717) begin
		AssumePrime = 1;
	end	else if (num==16'd32719) begin
		AssumePrime = 1;
	end	else if (num==16'd32749) begin
		AssumePrime = 1;
	end	else if (num==16'd32771) begin
		AssumePrime = 1;
	end	else if (num==16'd32779) begin
		AssumePrime = 1;
	end	else if (num==16'd32783) begin
		AssumePrime = 1;
	end	else if (num==16'd32789) begin
		AssumePrime = 1;
	end	else if (num==16'd32797) begin
		AssumePrime = 1;
	end	else if (num==16'd32801) begin
		AssumePrime = 1;
	end	else if (num==16'd32803) begin
		AssumePrime = 1;
	end	else if (num==16'd32831) begin
		AssumePrime = 1;
	end	else if (num==16'd32833) begin
		AssumePrime = 1;
	end	else if (num==16'd32839) begin
		AssumePrime = 1;
	end	else if (num==16'd32843) begin
		AssumePrime = 1;
	end	else if (num==16'd32869) begin
		AssumePrime = 1;
	end	else if (num==16'd32887) begin
		AssumePrime = 1;
	end	else if (num==16'd32909) begin
		AssumePrime = 1;
	end	else if (num==16'd32911) begin
		AssumePrime = 1;
	end	else if (num==16'd32917) begin
		AssumePrime = 1;
	end	else if (num==16'd32933) begin
		AssumePrime = 1;
	end	else if (num==16'd32939) begin
		AssumePrime = 1;
	end	else if (num==16'd32941) begin
		AssumePrime = 1;
	end	else if (num==16'd32957) begin
		AssumePrime = 1;
	end	else if (num==16'd32969) begin
		AssumePrime = 1;
	end	else if (num==16'd32971) begin
		AssumePrime = 1;
	end	else if (num==16'd32983) begin
		AssumePrime = 1;
	end	else if (num==16'd32987) begin
		AssumePrime = 1;
	end	else if (num==16'd32993) begin
		AssumePrime = 1;
	end	else if (num==16'd32999) begin
		AssumePrime = 1;
	end	else if (num==16'd33013) begin
		AssumePrime = 1;
	end	else if (num==16'd33023) begin
		AssumePrime = 1;
	end	else if (num==16'd33029) begin
		AssumePrime = 1;
	end	else if (num==16'd33037) begin
		AssumePrime = 1;
	end	else if (num==16'd33049) begin
		AssumePrime = 1;
	end	else if (num==16'd33053) begin
		AssumePrime = 1;
	end	else if (num==16'd33071) begin
		AssumePrime = 1;
	end	else if (num==16'd33073) begin
		AssumePrime = 1;
	end	else if (num==16'd33083) begin
		AssumePrime = 1;
	end	else if (num==16'd33091) begin
		AssumePrime = 1;
	end	else if (num==16'd33107) begin
		AssumePrime = 1;
	end	else if (num==16'd33113) begin
		AssumePrime = 1;
	end	else if (num==16'd33119) begin
		AssumePrime = 1;
	end	else if (num==16'd33149) begin
		AssumePrime = 1;
	end	else if (num==16'd33151) begin
		AssumePrime = 1;
	end	else if (num==16'd33161) begin
		AssumePrime = 1;
	end	else if (num==16'd33179) begin
		AssumePrime = 1;
	end	else if (num==16'd33181) begin
		AssumePrime = 1;
	end	else if (num==16'd33191) begin
		AssumePrime = 1;
	end	else if (num==16'd33199) begin
		AssumePrime = 1;
	end	else if (num==16'd33203) begin
		AssumePrime = 1;
	end	else if (num==16'd33211) begin
		AssumePrime = 1;
	end	else if (num==16'd33223) begin
		AssumePrime = 1;
	end	else if (num==16'd33247) begin
		AssumePrime = 1;
	end	else if (num==16'd33287) begin
		AssumePrime = 1;
	end	else if (num==16'd33289) begin
		AssumePrime = 1;
	end	else if (num==16'd33301) begin
		AssumePrime = 1;
	end	else if (num==16'd33311) begin
		AssumePrime = 1;
	end	else if (num==16'd33317) begin
		AssumePrime = 1;
	end	else if (num==16'd33329) begin
		AssumePrime = 1;
	end	else if (num==16'd33331) begin
		AssumePrime = 1;
	end	else if (num==16'd33343) begin
		AssumePrime = 1;
	end	else if (num==16'd33347) begin
		AssumePrime = 1;
	end	else if (num==16'd33349) begin
		AssumePrime = 1;
	end	else if (num==16'd33353) begin
		AssumePrime = 1;
	end	else if (num==16'd33359) begin
		AssumePrime = 1;
	end	else if (num==16'd33377) begin
		AssumePrime = 1;
	end	else if (num==16'd33391) begin
		AssumePrime = 1;
	end	else if (num==16'd33403) begin
		AssumePrime = 1;
	end	else if (num==16'd33409) begin
		AssumePrime = 1;
	end	else if (num==16'd33413) begin
		AssumePrime = 1;
	end	else if (num==16'd33427) begin
		AssumePrime = 1;
	end	else if (num==16'd33457) begin
		AssumePrime = 1;
	end	else if (num==16'd33461) begin
		AssumePrime = 1;
	end	else if (num==16'd33469) begin
		AssumePrime = 1;
	end	else if (num==16'd33479) begin
		AssumePrime = 1;
	end	else if (num==16'd33487) begin
		AssumePrime = 1;
	end	else if (num==16'd33493) begin
		AssumePrime = 1;
	end	else if (num==16'd33503) begin
		AssumePrime = 1;
	end	else if (num==16'd33521) begin
		AssumePrime = 1;
	end	else if (num==16'd33529) begin
		AssumePrime = 1;
	end	else if (num==16'd33533) begin
		AssumePrime = 1;
	end	else if (num==16'd33547) begin
		AssumePrime = 1;
	end	else if (num==16'd33563) begin
		AssumePrime = 1;
	end	else if (num==16'd33569) begin
		AssumePrime = 1;
	end	else if (num==16'd33577) begin
		AssumePrime = 1;
	end	else if (num==16'd33581) begin
		AssumePrime = 1;
	end	else if (num==16'd33587) begin
		AssumePrime = 1;
	end	else if (num==16'd33589) begin
		AssumePrime = 1;
	end	else if (num==16'd33599) begin
		AssumePrime = 1;
	end	else if (num==16'd33601) begin
		AssumePrime = 1;
	end	else if (num==16'd33613) begin
		AssumePrime = 1;
	end	else if (num==16'd33617) begin
		AssumePrime = 1;
	end	else if (num==16'd33619) begin
		AssumePrime = 1;
	end	else if (num==16'd33623) begin
		AssumePrime = 1;
	end	else if (num==16'd33629) begin
		AssumePrime = 1;
	end	else if (num==16'd33637) begin
		AssumePrime = 1;
	end	else if (num==16'd33641) begin
		AssumePrime = 1;
	end	else if (num==16'd33647) begin
		AssumePrime = 1;
	end	else if (num==16'd33679) begin
		AssumePrime = 1;
	end	else if (num==16'd33703) begin
		AssumePrime = 1;
	end	else if (num==16'd33713) begin
		AssumePrime = 1;
	end	else if (num==16'd33721) begin
		AssumePrime = 1;
	end	else if (num==16'd33739) begin
		AssumePrime = 1;
	end	else if (num==16'd33749) begin
		AssumePrime = 1;
	end	else if (num==16'd33751) begin
		AssumePrime = 1;
	end	else if (num==16'd33757) begin
		AssumePrime = 1;
	end	else if (num==16'd33767) begin
		AssumePrime = 1;
	end	else if (num==16'd33769) begin
		AssumePrime = 1;
	end	else if (num==16'd33773) begin
		AssumePrime = 1;
	end	else if (num==16'd33791) begin
		AssumePrime = 1;
	end	else if (num==16'd33797) begin
		AssumePrime = 1;
	end	else if (num==16'd33809) begin
		AssumePrime = 1;
	end	else if (num==16'd33811) begin
		AssumePrime = 1;
	end	else if (num==16'd33827) begin
		AssumePrime = 1;
	end	else if (num==16'd33829) begin
		AssumePrime = 1;
	end	else if (num==16'd33851) begin
		AssumePrime = 1;
	end	else if (num==16'd33857) begin
		AssumePrime = 1;
	end	else if (num==16'd33863) begin
		AssumePrime = 1;
	end	else if (num==16'd33871) begin
		AssumePrime = 1;
	end	else if (num==16'd33889) begin
		AssumePrime = 1;
	end	else if (num==16'd33893) begin
		AssumePrime = 1;
	end	else if (num==16'd33911) begin
		AssumePrime = 1;
	end	else if (num==16'd33923) begin
		AssumePrime = 1;
	end	else if (num==16'd33931) begin
		AssumePrime = 1;
	end	else if (num==16'd33937) begin
		AssumePrime = 1;
	end	else if (num==16'd33941) begin
		AssumePrime = 1;
	end	else if (num==16'd33961) begin
		AssumePrime = 1;
	end	else if (num==16'd33967) begin
		AssumePrime = 1;
	end	else if (num==16'd33997) begin
		AssumePrime = 1;
	end	else if (num==16'd34019) begin
		AssumePrime = 1;
	end	else if (num==16'd34031) begin
		AssumePrime = 1;
	end	else if (num==16'd34033) begin
		AssumePrime = 1;
	end	else if (num==16'd34039) begin
		AssumePrime = 1;
	end	else if (num==16'd34057) begin
		AssumePrime = 1;
	end	else if (num==16'd34061) begin
		AssumePrime = 1;
	end	else if (num==16'd34123) begin
		AssumePrime = 1;
	end	else if (num==16'd34127) begin
		AssumePrime = 1;
	end	else if (num==16'd34129) begin
		AssumePrime = 1;
	end	else if (num==16'd34141) begin
		AssumePrime = 1;
	end	else if (num==16'd34147) begin
		AssumePrime = 1;
	end	else if (num==16'd34157) begin
		AssumePrime = 1;
	end	else if (num==16'd34159) begin
		AssumePrime = 1;
	end	else if (num==16'd34171) begin
		AssumePrime = 1;
	end	else if (num==16'd34183) begin
		AssumePrime = 1;
	end	else if (num==16'd34211) begin
		AssumePrime = 1;
	end	else if (num==16'd34213) begin
		AssumePrime = 1;
	end	else if (num==16'd34217) begin
		AssumePrime = 1;
	end	else if (num==16'd34231) begin
		AssumePrime = 1;
	end	else if (num==16'd34253) begin
		AssumePrime = 1;
	end	else if (num==16'd34259) begin
		AssumePrime = 1;
	end	else if (num==16'd34261) begin
		AssumePrime = 1;
	end	else if (num==16'd34267) begin
		AssumePrime = 1;
	end	else if (num==16'd34273) begin
		AssumePrime = 1;
	end	else if (num==16'd34283) begin
		AssumePrime = 1;
	end	else if (num==16'd34297) begin
		AssumePrime = 1;
	end	else if (num==16'd34301) begin
		AssumePrime = 1;
	end	else if (num==16'd34303) begin
		AssumePrime = 1;
	end	else if (num==16'd34313) begin
		AssumePrime = 1;
	end	else if (num==16'd34319) begin
		AssumePrime = 1;
	end	else if (num==16'd34327) begin
		AssumePrime = 1;
	end	else if (num==16'd34337) begin
		AssumePrime = 1;
	end	else if (num==16'd34351) begin
		AssumePrime = 1;
	end	else if (num==16'd34361) begin
		AssumePrime = 1;
	end	else if (num==16'd34367) begin
		AssumePrime = 1;
	end	else if (num==16'd34369) begin
		AssumePrime = 1;
	end	else if (num==16'd34381) begin
		AssumePrime = 1;
	end	else if (num==16'd34403) begin
		AssumePrime = 1;
	end	else if (num==16'd34421) begin
		AssumePrime = 1;
	end	else if (num==16'd34429) begin
		AssumePrime = 1;
	end	else if (num==16'd34439) begin
		AssumePrime = 1;
	end	else if (num==16'd34457) begin
		AssumePrime = 1;
	end	else if (num==16'd34469) begin
		AssumePrime = 1;
	end	else if (num==16'd34471) begin
		AssumePrime = 1;
	end	else if (num==16'd34483) begin
		AssumePrime = 1;
	end	else if (num==16'd34487) begin
		AssumePrime = 1;
	end	else if (num==16'd34499) begin
		AssumePrime = 1;
	end	else if (num==16'd34501) begin
		AssumePrime = 1;
	end	else if (num==16'd34511) begin
		AssumePrime = 1;
	end	else if (num==16'd34513) begin
		AssumePrime = 1;
	end	else if (num==16'd34519) begin
		AssumePrime = 1;
	end	else if (num==16'd34537) begin
		AssumePrime = 1;
	end	else if (num==16'd34543) begin
		AssumePrime = 1;
	end	else if (num==16'd34549) begin
		AssumePrime = 1;
	end	else if (num==16'd34583) begin
		AssumePrime = 1;
	end	else if (num==16'd34589) begin
		AssumePrime = 1;
	end	else if (num==16'd34591) begin
		AssumePrime = 1;
	end	else if (num==16'd34603) begin
		AssumePrime = 1;
	end	else if (num==16'd34607) begin
		AssumePrime = 1;
	end	else if (num==16'd34613) begin
		AssumePrime = 1;
	end	else if (num==16'd34631) begin
		AssumePrime = 1;
	end	else if (num==16'd34649) begin
		AssumePrime = 1;
	end	else if (num==16'd34651) begin
		AssumePrime = 1;
	end	else if (num==16'd34667) begin
		AssumePrime = 1;
	end	else if (num==16'd34673) begin
		AssumePrime = 1;
	end	else if (num==16'd34679) begin
		AssumePrime = 1;
	end	else if (num==16'd34687) begin
		AssumePrime = 1;
	end	else if (num==16'd34693) begin
		AssumePrime = 1;
	end	else if (num==16'd34703) begin
		AssumePrime = 1;
	end	else if (num==16'd34721) begin
		AssumePrime = 1;
	end	else if (num==16'd34729) begin
		AssumePrime = 1;
	end	else if (num==16'd34739) begin
		AssumePrime = 1;
	end	else if (num==16'd34747) begin
		AssumePrime = 1;
	end	else if (num==16'd34757) begin
		AssumePrime = 1;
	end	else if (num==16'd34759) begin
		AssumePrime = 1;
	end	else if (num==16'd34763) begin
		AssumePrime = 1;
	end	else if (num==16'd34781) begin
		AssumePrime = 1;
	end	else if (num==16'd34807) begin
		AssumePrime = 1;
	end	else if (num==16'd34819) begin
		AssumePrime = 1;
	end	else if (num==16'd34841) begin
		AssumePrime = 1;
	end	else if (num==16'd34843) begin
		AssumePrime = 1;
	end	else if (num==16'd34847) begin
		AssumePrime = 1;
	end	else if (num==16'd34849) begin
		AssumePrime = 1;
	end	else if (num==16'd34871) begin
		AssumePrime = 1;
	end	else if (num==16'd34877) begin
		AssumePrime = 1;
	end	else if (num==16'd34883) begin
		AssumePrime = 1;
	end	else if (num==16'd34897) begin
		AssumePrime = 1;
	end	else if (num==16'd34913) begin
		AssumePrime = 1;
	end	else if (num==16'd34919) begin
		AssumePrime = 1;
	end	else if (num==16'd34939) begin
		AssumePrime = 1;
	end	else if (num==16'd34949) begin
		AssumePrime = 1;
	end	else if (num==16'd34961) begin
		AssumePrime = 1;
	end	else if (num==16'd34963) begin
		AssumePrime = 1;
	end	else if (num==16'd34981) begin
		AssumePrime = 1;
	end	else if (num==16'd35023) begin
		AssumePrime = 1;
	end	else if (num==16'd35027) begin
		AssumePrime = 1;
	end	else if (num==16'd35051) begin
		AssumePrime = 1;
	end	else if (num==16'd35053) begin
		AssumePrime = 1;
	end	else if (num==16'd35059) begin
		AssumePrime = 1;
	end	else if (num==16'd35069) begin
		AssumePrime = 1;
	end	else if (num==16'd35081) begin
		AssumePrime = 1;
	end	else if (num==16'd35083) begin
		AssumePrime = 1;
	end	else if (num==16'd35089) begin
		AssumePrime = 1;
	end	else if (num==16'd35099) begin
		AssumePrime = 1;
	end	else if (num==16'd35107) begin
		AssumePrime = 1;
	end	else if (num==16'd35111) begin
		AssumePrime = 1;
	end	else if (num==16'd35117) begin
		AssumePrime = 1;
	end	else if (num==16'd35129) begin
		AssumePrime = 1;
	end	else if (num==16'd35141) begin
		AssumePrime = 1;
	end	else if (num==16'd35149) begin
		AssumePrime = 1;
	end	else if (num==16'd35153) begin
		AssumePrime = 1;
	end	else if (num==16'd35159) begin
		AssumePrime = 1;
	end	else if (num==16'd35171) begin
		AssumePrime = 1;
	end	else if (num==16'd35201) begin
		AssumePrime = 1;
	end	else if (num==16'd35221) begin
		AssumePrime = 1;
	end	else if (num==16'd35227) begin
		AssumePrime = 1;
	end	else if (num==16'd35251) begin
		AssumePrime = 1;
	end	else if (num==16'd35257) begin
		AssumePrime = 1;
	end	else if (num==16'd35267) begin
		AssumePrime = 1;
	end	else if (num==16'd35279) begin
		AssumePrime = 1;
	end	else if (num==16'd35281) begin
		AssumePrime = 1;
	end	else if (num==16'd35291) begin
		AssumePrime = 1;
	end	else if (num==16'd35311) begin
		AssumePrime = 1;
	end	else if (num==16'd35317) begin
		AssumePrime = 1;
	end	else if (num==16'd35323) begin
		AssumePrime = 1;
	end	else if (num==16'd35327) begin
		AssumePrime = 1;
	end	else if (num==16'd35339) begin
		AssumePrime = 1;
	end	else if (num==16'd35353) begin
		AssumePrime = 1;
	end	else if (num==16'd35363) begin
		AssumePrime = 1;
	end	else if (num==16'd35381) begin
		AssumePrime = 1;
	end	else if (num==16'd35393) begin
		AssumePrime = 1;
	end	else if (num==16'd35401) begin
		AssumePrime = 1;
	end	else if (num==16'd35407) begin
		AssumePrime = 1;
	end	else if (num==16'd35419) begin
		AssumePrime = 1;
	end	else if (num==16'd35423) begin
		AssumePrime = 1;
	end	else if (num==16'd35437) begin
		AssumePrime = 1;
	end	else if (num==16'd35447) begin
		AssumePrime = 1;
	end	else if (num==16'd35449) begin
		AssumePrime = 1;
	end	else if (num==16'd35461) begin
		AssumePrime = 1;
	end	else if (num==16'd35491) begin
		AssumePrime = 1;
	end	else if (num==16'd35507) begin
		AssumePrime = 1;
	end	else if (num==16'd35509) begin
		AssumePrime = 1;
	end	else if (num==16'd35521) begin
		AssumePrime = 1;
	end	else if (num==16'd35527) begin
		AssumePrime = 1;
	end	else if (num==16'd35531) begin
		AssumePrime = 1;
	end	else if (num==16'd35533) begin
		AssumePrime = 1;
	end	else if (num==16'd35537) begin
		AssumePrime = 1;
	end	else if (num==16'd35543) begin
		AssumePrime = 1;
	end	else if (num==16'd35569) begin
		AssumePrime = 1;
	end	else if (num==16'd35573) begin
		AssumePrime = 1;
	end	else if (num==16'd35591) begin
		AssumePrime = 1;
	end	else if (num==16'd35593) begin
		AssumePrime = 1;
	end	else if (num==16'd35597) begin
		AssumePrime = 1;
	end	else if (num==16'd35603) begin
		AssumePrime = 1;
	end	else if (num==16'd35617) begin
		AssumePrime = 1;
	end	else if (num==16'd35671) begin
		AssumePrime = 1;
	end	else if (num==16'd35677) begin
		AssumePrime = 1;
	end	else if (num==16'd35729) begin
		AssumePrime = 1;
	end	else if (num==16'd35731) begin
		AssumePrime = 1;
	end	else if (num==16'd35747) begin
		AssumePrime = 1;
	end	else if (num==16'd35753) begin
		AssumePrime = 1;
	end	else if (num==16'd35759) begin
		AssumePrime = 1;
	end	else if (num==16'd35771) begin
		AssumePrime = 1;
	end	else if (num==16'd35797) begin
		AssumePrime = 1;
	end	else if (num==16'd35801) begin
		AssumePrime = 1;
	end	else if (num==16'd35803) begin
		AssumePrime = 1;
	end	else if (num==16'd35809) begin
		AssumePrime = 1;
	end	else if (num==16'd35831) begin
		AssumePrime = 1;
	end	else if (num==16'd35837) begin
		AssumePrime = 1;
	end	else if (num==16'd35839) begin
		AssumePrime = 1;
	end	else if (num==16'd35851) begin
		AssumePrime = 1;
	end	else if (num==16'd35863) begin
		AssumePrime = 1;
	end	else if (num==16'd35869) begin
		AssumePrime = 1;
	end	else if (num==16'd35879) begin
		AssumePrime = 1;
	end	else if (num==16'd35897) begin
		AssumePrime = 1;
	end	else if (num==16'd35899) begin
		AssumePrime = 1;
	end	else if (num==16'd35911) begin
		AssumePrime = 1;
	end	else if (num==16'd35923) begin
		AssumePrime = 1;
	end	else if (num==16'd35933) begin
		AssumePrime = 1;
	end	else if (num==16'd35951) begin
		AssumePrime = 1;
	end	else if (num==16'd35963) begin
		AssumePrime = 1;
	end	else if (num==16'd35969) begin
		AssumePrime = 1;
	end	else if (num==16'd35977) begin
		AssumePrime = 1;
	end	else if (num==16'd35983) begin
		AssumePrime = 1;
	end	else if (num==16'd35993) begin
		AssumePrime = 1;
	end	else if (num==16'd35999) begin
		AssumePrime = 1;
	end	else if (num==16'd36007) begin
		AssumePrime = 1;
	end	else if (num==16'd36011) begin
		AssumePrime = 1;
	end	else if (num==16'd36013) begin
		AssumePrime = 1;
	end	else if (num==16'd36017) begin
		AssumePrime = 1;
	end	else if (num==16'd36037) begin
		AssumePrime = 1;
	end	else if (num==16'd36061) begin
		AssumePrime = 1;
	end	else if (num==16'd36067) begin
		AssumePrime = 1;
	end	else if (num==16'd36073) begin
		AssumePrime = 1;
	end	else if (num==16'd36083) begin
		AssumePrime = 1;
	end	else if (num==16'd36097) begin
		AssumePrime = 1;
	end	else if (num==16'd36107) begin
		AssumePrime = 1;
	end	else if (num==16'd36109) begin
		AssumePrime = 1;
	end	else if (num==16'd36131) begin
		AssumePrime = 1;
	end	else if (num==16'd36137) begin
		AssumePrime = 1;
	end	else if (num==16'd36151) begin
		AssumePrime = 1;
	end	else if (num==16'd36161) begin
		AssumePrime = 1;
	end	else if (num==16'd36187) begin
		AssumePrime = 1;
	end	else if (num==16'd36191) begin
		AssumePrime = 1;
	end	else if (num==16'd36209) begin
		AssumePrime = 1;
	end	else if (num==16'd36217) begin
		AssumePrime = 1;
	end	else if (num==16'd36229) begin
		AssumePrime = 1;
	end	else if (num==16'd36241) begin
		AssumePrime = 1;
	end	else if (num==16'd36251) begin
		AssumePrime = 1;
	end	else if (num==16'd36263) begin
		AssumePrime = 1;
	end	else if (num==16'd36269) begin
		AssumePrime = 1;
	end	else if (num==16'd36277) begin
		AssumePrime = 1;
	end	else if (num==16'd36293) begin
		AssumePrime = 1;
	end	else if (num==16'd36299) begin
		AssumePrime = 1;
	end	else if (num==16'd36307) begin
		AssumePrime = 1;
	end	else if (num==16'd36313) begin
		AssumePrime = 1;
	end	else if (num==16'd36319) begin
		AssumePrime = 1;
	end	else if (num==16'd36341) begin
		AssumePrime = 1;
	end	else if (num==16'd36343) begin
		AssumePrime = 1;
	end	else if (num==16'd36353) begin
		AssumePrime = 1;
	end	else if (num==16'd36373) begin
		AssumePrime = 1;
	end	else if (num==16'd36383) begin
		AssumePrime = 1;
	end	else if (num==16'd36389) begin
		AssumePrime = 1;
	end	else if (num==16'd36433) begin
		AssumePrime = 1;
	end	else if (num==16'd36451) begin
		AssumePrime = 1;
	end	else if (num==16'd36457) begin
		AssumePrime = 1;
	end	else if (num==16'd36467) begin
		AssumePrime = 1;
	end	else if (num==16'd36469) begin
		AssumePrime = 1;
	end	else if (num==16'd36473) begin
		AssumePrime = 1;
	end	else if (num==16'd36479) begin
		AssumePrime = 1;
	end	else if (num==16'd36493) begin
		AssumePrime = 1;
	end	else if (num==16'd36497) begin
		AssumePrime = 1;
	end	else if (num==16'd36523) begin
		AssumePrime = 1;
	end	else if (num==16'd36527) begin
		AssumePrime = 1;
	end	else if (num==16'd36529) begin
		AssumePrime = 1;
	end	else if (num==16'd36541) begin
		AssumePrime = 1;
	end	else if (num==16'd36551) begin
		AssumePrime = 1;
	end	else if (num==16'd36559) begin
		AssumePrime = 1;
	end	else if (num==16'd36563) begin
		AssumePrime = 1;
	end	else if (num==16'd36571) begin
		AssumePrime = 1;
	end	else if (num==16'd36583) begin
		AssumePrime = 1;
	end	else if (num==16'd36587) begin
		AssumePrime = 1;
	end	else if (num==16'd36599) begin
		AssumePrime = 1;
	end	else if (num==16'd36607) begin
		AssumePrime = 1;
	end	else if (num==16'd36629) begin
		AssumePrime = 1;
	end	else if (num==16'd36637) begin
		AssumePrime = 1;
	end	else if (num==16'd36643) begin
		AssumePrime = 1;
	end	else if (num==16'd36653) begin
		AssumePrime = 1;
	end	else if (num==16'd36671) begin
		AssumePrime = 1;
	end	else if (num==16'd36677) begin
		AssumePrime = 1;
	end	else if (num==16'd36683) begin
		AssumePrime = 1;
	end	else if (num==16'd36691) begin
		AssumePrime = 1;
	end	else if (num==16'd36697) begin
		AssumePrime = 1;
	end	else if (num==16'd36709) begin
		AssumePrime = 1;
	end	else if (num==16'd36713) begin
		AssumePrime = 1;
	end	else if (num==16'd36721) begin
		AssumePrime = 1;
	end	else if (num==16'd36739) begin
		AssumePrime = 1;
	end	else if (num==16'd36749) begin
		AssumePrime = 1;
	end	else if (num==16'd36761) begin
		AssumePrime = 1;
	end	else if (num==16'd36767) begin
		AssumePrime = 1;
	end	else if (num==16'd36779) begin
		AssumePrime = 1;
	end	else if (num==16'd36781) begin
		AssumePrime = 1;
	end	else if (num==16'd36787) begin
		AssumePrime = 1;
	end	else if (num==16'd36791) begin
		AssumePrime = 1;
	end	else if (num==16'd36793) begin
		AssumePrime = 1;
	end	else if (num==16'd36809) begin
		AssumePrime = 1;
	end	else if (num==16'd36821) begin
		AssumePrime = 1;
	end	else if (num==16'd36833) begin
		AssumePrime = 1;
	end	else if (num==16'd36847) begin
		AssumePrime = 1;
	end	else if (num==16'd36857) begin
		AssumePrime = 1;
	end	else if (num==16'd36871) begin
		AssumePrime = 1;
	end	else if (num==16'd36877) begin
		AssumePrime = 1;
	end	else if (num==16'd36887) begin
		AssumePrime = 1;
	end	else if (num==16'd36899) begin
		AssumePrime = 1;
	end	else if (num==16'd36901) begin
		AssumePrime = 1;
	end	else if (num==16'd36913) begin
		AssumePrime = 1;
	end	else if (num==16'd36919) begin
		AssumePrime = 1;
	end	else if (num==16'd36923) begin
		AssumePrime = 1;
	end	else if (num==16'd36929) begin
		AssumePrime = 1;
	end	else if (num==16'd36931) begin
		AssumePrime = 1;
	end	else if (num==16'd36943) begin
		AssumePrime = 1;
	end	else if (num==16'd36947) begin
		AssumePrime = 1;
	end	else if (num==16'd36973) begin
		AssumePrime = 1;
	end	else if (num==16'd36979) begin
		AssumePrime = 1;
	end	else if (num==16'd36997) begin
		AssumePrime = 1;
	end	else if (num==16'd37003) begin
		AssumePrime = 1;
	end	else if (num==16'd37013) begin
		AssumePrime = 1;
	end	else if (num==16'd37019) begin
		AssumePrime = 1;
	end	else if (num==16'd37021) begin
		AssumePrime = 1;
	end	else if (num==16'd37039) begin
		AssumePrime = 1;
	end	else if (num==16'd37049) begin
		AssumePrime = 1;
	end	else if (num==16'd37057) begin
		AssumePrime = 1;
	end	else if (num==16'd37061) begin
		AssumePrime = 1;
	end	else if (num==16'd37087) begin
		AssumePrime = 1;
	end	else if (num==16'd37097) begin
		AssumePrime = 1;
	end	else if (num==16'd37117) begin
		AssumePrime = 1;
	end	else if (num==16'd37123) begin
		AssumePrime = 1;
	end	else if (num==16'd37139) begin
		AssumePrime = 1;
	end	else if (num==16'd37159) begin
		AssumePrime = 1;
	end	else if (num==16'd37171) begin
		AssumePrime = 1;
	end	else if (num==16'd37181) begin
		AssumePrime = 1;
	end	else if (num==16'd37189) begin
		AssumePrime = 1;
	end	else if (num==16'd37199) begin
		AssumePrime = 1;
	end	else if (num==16'd37201) begin
		AssumePrime = 1;
	end	else if (num==16'd37217) begin
		AssumePrime = 1;
	end	else if (num==16'd37223) begin
		AssumePrime = 1;
	end	else if (num==16'd37243) begin
		AssumePrime = 1;
	end	else if (num==16'd37253) begin
		AssumePrime = 1;
	end	else if (num==16'd37273) begin
		AssumePrime = 1;
	end	else if (num==16'd37277) begin
		AssumePrime = 1;
	end	else if (num==16'd37307) begin
		AssumePrime = 1;
	end	else if (num==16'd37309) begin
		AssumePrime = 1;
	end	else if (num==16'd37313) begin
		AssumePrime = 1;
	end	else if (num==16'd37321) begin
		AssumePrime = 1;
	end	else if (num==16'd37337) begin
		AssumePrime = 1;
	end	else if (num==16'd37339) begin
		AssumePrime = 1;
	end	else if (num==16'd37357) begin
		AssumePrime = 1;
	end	else if (num==16'd37361) begin
		AssumePrime = 1;
	end	else if (num==16'd37363) begin
		AssumePrime = 1;
	end	else if (num==16'd37369) begin
		AssumePrime = 1;
	end	else if (num==16'd37379) begin
		AssumePrime = 1;
	end	else if (num==16'd37397) begin
		AssumePrime = 1;
	end	else if (num==16'd37409) begin
		AssumePrime = 1;
	end	else if (num==16'd37423) begin
		AssumePrime = 1;
	end	else if (num==16'd37441) begin
		AssumePrime = 1;
	end	else if (num==16'd37447) begin
		AssumePrime = 1;
	end	else if (num==16'd37463) begin
		AssumePrime = 1;
	end	else if (num==16'd37483) begin
		AssumePrime = 1;
	end	else if (num==16'd37489) begin
		AssumePrime = 1;
	end	else if (num==16'd37493) begin
		AssumePrime = 1;
	end	else if (num==16'd37501) begin
		AssumePrime = 1;
	end	else if (num==16'd37507) begin
		AssumePrime = 1;
	end	else if (num==16'd37511) begin
		AssumePrime = 1;
	end	else if (num==16'd37517) begin
		AssumePrime = 1;
	end	else if (num==16'd37529) begin
		AssumePrime = 1;
	end	else if (num==16'd37537) begin
		AssumePrime = 1;
	end	else if (num==16'd37547) begin
		AssumePrime = 1;
	end	else if (num==16'd37549) begin
		AssumePrime = 1;
	end	else if (num==16'd37561) begin
		AssumePrime = 1;
	end	else if (num==16'd37567) begin
		AssumePrime = 1;
	end	else if (num==16'd37571) begin
		AssumePrime = 1;
	end	else if (num==16'd37573) begin
		AssumePrime = 1;
	end	else if (num==16'd37579) begin
		AssumePrime = 1;
	end	else if (num==16'd37589) begin
		AssumePrime = 1;
	end	else if (num==16'd37591) begin
		AssumePrime = 1;
	end	else if (num==16'd37607) begin
		AssumePrime = 1;
	end	else if (num==16'd37619) begin
		AssumePrime = 1;
	end	else if (num==16'd37633) begin
		AssumePrime = 1;
	end	else if (num==16'd37643) begin
		AssumePrime = 1;
	end	else if (num==16'd37649) begin
		AssumePrime = 1;
	end	else if (num==16'd37657) begin
		AssumePrime = 1;
	end	else if (num==16'd37663) begin
		AssumePrime = 1;
	end	else if (num==16'd37691) begin
		AssumePrime = 1;
	end	else if (num==16'd37693) begin
		AssumePrime = 1;
	end	else if (num==16'd37699) begin
		AssumePrime = 1;
	end	else if (num==16'd37717) begin
		AssumePrime = 1;
	end	else if (num==16'd37747) begin
		AssumePrime = 1;
	end	else if (num==16'd37781) begin
		AssumePrime = 1;
	end	else if (num==16'd37783) begin
		AssumePrime = 1;
	end	else if (num==16'd37799) begin
		AssumePrime = 1;
	end	else if (num==16'd37811) begin
		AssumePrime = 1;
	end	else if (num==16'd37813) begin
		AssumePrime = 1;
	end	else if (num==16'd37831) begin
		AssumePrime = 1;
	end	else if (num==16'd37847) begin
		AssumePrime = 1;
	end	else if (num==16'd37853) begin
		AssumePrime = 1;
	end	else if (num==16'd37861) begin
		AssumePrime = 1;
	end	else if (num==16'd37871) begin
		AssumePrime = 1;
	end	else if (num==16'd37879) begin
		AssumePrime = 1;
	end	else if (num==16'd37889) begin
		AssumePrime = 1;
	end	else if (num==16'd37897) begin
		AssumePrime = 1;
	end	else if (num==16'd37907) begin
		AssumePrime = 1;
	end	else if (num==16'd37951) begin
		AssumePrime = 1;
	end	else if (num==16'd37957) begin
		AssumePrime = 1;
	end	else if (num==16'd37963) begin
		AssumePrime = 1;
	end	else if (num==16'd37967) begin
		AssumePrime = 1;
	end	else if (num==16'd37987) begin
		AssumePrime = 1;
	end	else if (num==16'd37991) begin
		AssumePrime = 1;
	end	else if (num==16'd37993) begin
		AssumePrime = 1;
	end	else if (num==16'd37997) begin
		AssumePrime = 1;
	end	else if (num==16'd38011) begin
		AssumePrime = 1;
	end	else if (num==16'd38039) begin
		AssumePrime = 1;
	end	else if (num==16'd38047) begin
		AssumePrime = 1;
	end	else if (num==16'd38053) begin
		AssumePrime = 1;
	end	else if (num==16'd38069) begin
		AssumePrime = 1;
	end	else if (num==16'd38083) begin
		AssumePrime = 1;
	end	else if (num==16'd38113) begin
		AssumePrime = 1;
	end	else if (num==16'd38119) begin
		AssumePrime = 1;
	end	else if (num==16'd38149) begin
		AssumePrime = 1;
	end	else if (num==16'd38153) begin
		AssumePrime = 1;
	end	else if (num==16'd38167) begin
		AssumePrime = 1;
	end	else if (num==16'd38177) begin
		AssumePrime = 1;
	end	else if (num==16'd38183) begin
		AssumePrime = 1;
	end	else if (num==16'd38189) begin
		AssumePrime = 1;
	end	else if (num==16'd38197) begin
		AssumePrime = 1;
	end	else if (num==16'd38201) begin
		AssumePrime = 1;
	end	else if (num==16'd38219) begin
		AssumePrime = 1;
	end	else if (num==16'd38231) begin
		AssumePrime = 1;
	end	else if (num==16'd38237) begin
		AssumePrime = 1;
	end	else if (num==16'd38239) begin
		AssumePrime = 1;
	end	else if (num==16'd38261) begin
		AssumePrime = 1;
	end	else if (num==16'd38273) begin
		AssumePrime = 1;
	end	else if (num==16'd38281) begin
		AssumePrime = 1;
	end	else if (num==16'd38287) begin
		AssumePrime = 1;
	end	else if (num==16'd38299) begin
		AssumePrime = 1;
	end	else if (num==16'd38303) begin
		AssumePrime = 1;
	end	else if (num==16'd38317) begin
		AssumePrime = 1;
	end	else if (num==16'd38321) begin
		AssumePrime = 1;
	end	else if (num==16'd38327) begin
		AssumePrime = 1;
	end	else if (num==16'd38329) begin
		AssumePrime = 1;
	end	else if (num==16'd38333) begin
		AssumePrime = 1;
	end	else if (num==16'd38351) begin
		AssumePrime = 1;
	end	else if (num==16'd38371) begin
		AssumePrime = 1;
	end	else if (num==16'd38377) begin
		AssumePrime = 1;
	end	else if (num==16'd38393) begin
		AssumePrime = 1;
	end	else if (num==16'd38431) begin
		AssumePrime = 1;
	end	else if (num==16'd38447) begin
		AssumePrime = 1;
	end	else if (num==16'd38449) begin
		AssumePrime = 1;
	end	else if (num==16'd38453) begin
		AssumePrime = 1;
	end	else if (num==16'd38459) begin
		AssumePrime = 1;
	end	else if (num==16'd38461) begin
		AssumePrime = 1;
	end	else if (num==16'd38501) begin
		AssumePrime = 1;
	end	else if (num==16'd38543) begin
		AssumePrime = 1;
	end	else if (num==16'd38557) begin
		AssumePrime = 1;
	end	else if (num==16'd38561) begin
		AssumePrime = 1;
	end	else if (num==16'd38567) begin
		AssumePrime = 1;
	end	else if (num==16'd38569) begin
		AssumePrime = 1;
	end	else if (num==16'd38593) begin
		AssumePrime = 1;
	end	else if (num==16'd38603) begin
		AssumePrime = 1;
	end	else if (num==16'd38609) begin
		AssumePrime = 1;
	end	else if (num==16'd38611) begin
		AssumePrime = 1;
	end	else if (num==16'd38629) begin
		AssumePrime = 1;
	end	else if (num==16'd38639) begin
		AssumePrime = 1;
	end	else if (num==16'd38651) begin
		AssumePrime = 1;
	end	else if (num==16'd38653) begin
		AssumePrime = 1;
	end	else if (num==16'd38669) begin
		AssumePrime = 1;
	end	else if (num==16'd38671) begin
		AssumePrime = 1;
	end	else if (num==16'd38677) begin
		AssumePrime = 1;
	end	else if (num==16'd38693) begin
		AssumePrime = 1;
	end	else if (num==16'd38699) begin
		AssumePrime = 1;
	end	else if (num==16'd38707) begin
		AssumePrime = 1;
	end	else if (num==16'd38711) begin
		AssumePrime = 1;
	end	else if (num==16'd38713) begin
		AssumePrime = 1;
	end	else if (num==16'd38723) begin
		AssumePrime = 1;
	end	else if (num==16'd38729) begin
		AssumePrime = 1;
	end	else if (num==16'd38737) begin
		AssumePrime = 1;
	end	else if (num==16'd38747) begin
		AssumePrime = 1;
	end	else if (num==16'd38749) begin
		AssumePrime = 1;
	end	else if (num==16'd38767) begin
		AssumePrime = 1;
	end	else if (num==16'd38783) begin
		AssumePrime = 1;
	end	else if (num==16'd38791) begin
		AssumePrime = 1;
	end	else if (num==16'd38803) begin
		AssumePrime = 1;
	end	else if (num==16'd38821) begin
		AssumePrime = 1;
	end	else if (num==16'd38833) begin
		AssumePrime = 1;
	end	else if (num==16'd38839) begin
		AssumePrime = 1;
	end	else if (num==16'd38851) begin
		AssumePrime = 1;
	end	else if (num==16'd38861) begin
		AssumePrime = 1;
	end	else if (num==16'd38867) begin
		AssumePrime = 1;
	end	else if (num==16'd38873) begin
		AssumePrime = 1;
	end	else if (num==16'd38891) begin
		AssumePrime = 1;
	end	else if (num==16'd38903) begin
		AssumePrime = 1;
	end	else if (num==16'd38917) begin
		AssumePrime = 1;
	end	else if (num==16'd38921) begin
		AssumePrime = 1;
	end	else if (num==16'd38923) begin
		AssumePrime = 1;
	end	else if (num==16'd38933) begin
		AssumePrime = 1;
	end	else if (num==16'd38953) begin
		AssumePrime = 1;
	end	else if (num==16'd38959) begin
		AssumePrime = 1;
	end	else if (num==16'd38971) begin
		AssumePrime = 1;
	end	else if (num==16'd38977) begin
		AssumePrime = 1;
	end	else if (num==16'd38993) begin
		AssumePrime = 1;
	end	else if (num==16'd39019) begin
		AssumePrime = 1;
	end	else if (num==16'd39023) begin
		AssumePrime = 1;
	end	else if (num==16'd39041) begin
		AssumePrime = 1;
	end	else if (num==16'd39043) begin
		AssumePrime = 1;
	end	else if (num==16'd39047) begin
		AssumePrime = 1;
	end	else if (num==16'd39079) begin
		AssumePrime = 1;
	end	else if (num==16'd39089) begin
		AssumePrime = 1;
	end	else if (num==16'd39097) begin
		AssumePrime = 1;
	end	else if (num==16'd39103) begin
		AssumePrime = 1;
	end	else if (num==16'd39107) begin
		AssumePrime = 1;
	end	else if (num==16'd39113) begin
		AssumePrime = 1;
	end	else if (num==16'd39119) begin
		AssumePrime = 1;
	end	else if (num==16'd39133) begin
		AssumePrime = 1;
	end	else if (num==16'd39139) begin
		AssumePrime = 1;
	end	else if (num==16'd39157) begin
		AssumePrime = 1;
	end	else if (num==16'd39161) begin
		AssumePrime = 1;
	end	else if (num==16'd39163) begin
		AssumePrime = 1;
	end	else if (num==16'd39181) begin
		AssumePrime = 1;
	end	else if (num==16'd39191) begin
		AssumePrime = 1;
	end	else if (num==16'd39199) begin
		AssumePrime = 1;
	end	else if (num==16'd39209) begin
		AssumePrime = 1;
	end	else if (num==16'd39217) begin
		AssumePrime = 1;
	end	else if (num==16'd39227) begin
		AssumePrime = 1;
	end	else if (num==16'd39229) begin
		AssumePrime = 1;
	end	else if (num==16'd39233) begin
		AssumePrime = 1;
	end	else if (num==16'd39239) begin
		AssumePrime = 1;
	end	else if (num==16'd39241) begin
		AssumePrime = 1;
	end	else if (num==16'd39251) begin
		AssumePrime = 1;
	end	else if (num==16'd39293) begin
		AssumePrime = 1;
	end	else if (num==16'd39301) begin
		AssumePrime = 1;
	end	else if (num==16'd39313) begin
		AssumePrime = 1;
	end	else if (num==16'd39317) begin
		AssumePrime = 1;
	end	else if (num==16'd39323) begin
		AssumePrime = 1;
	end	else if (num==16'd39341) begin
		AssumePrime = 1;
	end	else if (num==16'd39343) begin
		AssumePrime = 1;
	end	else if (num==16'd39359) begin
		AssumePrime = 1;
	end	else if (num==16'd39367) begin
		AssumePrime = 1;
	end	else if (num==16'd39371) begin
		AssumePrime = 1;
	end	else if (num==16'd39373) begin
		AssumePrime = 1;
	end	else if (num==16'd39383) begin
		AssumePrime = 1;
	end	else if (num==16'd39397) begin
		AssumePrime = 1;
	end	else if (num==16'd39409) begin
		AssumePrime = 1;
	end	else if (num==16'd39419) begin
		AssumePrime = 1;
	end	else if (num==16'd39439) begin
		AssumePrime = 1;
	end	else if (num==16'd39443) begin
		AssumePrime = 1;
	end	else if (num==16'd39451) begin
		AssumePrime = 1;
	end	else if (num==16'd39461) begin
		AssumePrime = 1;
	end	else if (num==16'd39499) begin
		AssumePrime = 1;
	end	else if (num==16'd39503) begin
		AssumePrime = 1;
	end	else if (num==16'd39509) begin
		AssumePrime = 1;
	end	else if (num==16'd39511) begin
		AssumePrime = 1;
	end	else if (num==16'd39521) begin
		AssumePrime = 1;
	end	else if (num==16'd39541) begin
		AssumePrime = 1;
	end	else if (num==16'd39551) begin
		AssumePrime = 1;
	end	else if (num==16'd39563) begin
		AssumePrime = 1;
	end	else if (num==16'd39569) begin
		AssumePrime = 1;
	end	else if (num==16'd39581) begin
		AssumePrime = 1;
	end	else if (num==16'd39607) begin
		AssumePrime = 1;
	end	else if (num==16'd39619) begin
		AssumePrime = 1;
	end	else if (num==16'd39623) begin
		AssumePrime = 1;
	end	else if (num==16'd39631) begin
		AssumePrime = 1;
	end	else if (num==16'd39659) begin
		AssumePrime = 1;
	end	else if (num==16'd39667) begin
		AssumePrime = 1;
	end	else if (num==16'd39671) begin
		AssumePrime = 1;
	end	else if (num==16'd39679) begin
		AssumePrime = 1;
	end	else if (num==16'd39703) begin
		AssumePrime = 1;
	end	else if (num==16'd39709) begin
		AssumePrime = 1;
	end	else if (num==16'd39719) begin
		AssumePrime = 1;
	end	else if (num==16'd39727) begin
		AssumePrime = 1;
	end	else if (num==16'd39733) begin
		AssumePrime = 1;
	end	else if (num==16'd39749) begin
		AssumePrime = 1;
	end	else if (num==16'd39761) begin
		AssumePrime = 1;
	end	else if (num==16'd39769) begin
		AssumePrime = 1;
	end	else if (num==16'd39779) begin
		AssumePrime = 1;
	end	else if (num==16'd39791) begin
		AssumePrime = 1;
	end	else if (num==16'd39799) begin
		AssumePrime = 1;
	end	else if (num==16'd39821) begin
		AssumePrime = 1;
	end	else if (num==16'd39827) begin
		AssumePrime = 1;
	end	else if (num==16'd39829) begin
		AssumePrime = 1;
	end	else if (num==16'd39839) begin
		AssumePrime = 1;
	end	else if (num==16'd39841) begin
		AssumePrime = 1;
	end	else if (num==16'd39847) begin
		AssumePrime = 1;
	end	else if (num==16'd39857) begin
		AssumePrime = 1;
	end	else if (num==16'd39863) begin
		AssumePrime = 1;
	end	else if (num==16'd39869) begin
		AssumePrime = 1;
	end	else if (num==16'd39877) begin
		AssumePrime = 1;
	end	else if (num==16'd39883) begin
		AssumePrime = 1;
	end	else if (num==16'd39887) begin
		AssumePrime = 1;
	end	else if (num==16'd39901) begin
		AssumePrime = 1;
	end	else if (num==16'd39929) begin
		AssumePrime = 1;
	end	else if (num==16'd39937) begin
		AssumePrime = 1;
	end	else if (num==16'd39953) begin
		AssumePrime = 1;
	end	else if (num==16'd39971) begin
		AssumePrime = 1;
	end	else if (num==16'd39979) begin
		AssumePrime = 1;
	end	else if (num==16'd39983) begin
		AssumePrime = 1;
	end	else if (num==16'd39989) begin
		AssumePrime = 1;
	end	else if (num==16'd40009) begin
		AssumePrime = 1;
	end	else if (num==16'd40013) begin
		AssumePrime = 1;
	end	else if (num==16'd40031) begin
		AssumePrime = 1;
	end	else if (num==16'd40037) begin
		AssumePrime = 1;
	end	else if (num==16'd40039) begin
		AssumePrime = 1;
	end	else if (num==16'd40063) begin
		AssumePrime = 1;
	end	else if (num==16'd40087) begin
		AssumePrime = 1;
	end	else if (num==16'd40093) begin
		AssumePrime = 1;
	end	else if (num==16'd40099) begin
		AssumePrime = 1;
	end	else if (num==16'd40111) begin
		AssumePrime = 1;
	end	else if (num==16'd40123) begin
		AssumePrime = 1;
	end	else if (num==16'd40127) begin
		AssumePrime = 1;
	end	else if (num==16'd40129) begin
		AssumePrime = 1;
	end	else if (num==16'd40151) begin
		AssumePrime = 1;
	end	else if (num==16'd40153) begin
		AssumePrime = 1;
	end	else if (num==16'd40163) begin
		AssumePrime = 1;
	end	else if (num==16'd40169) begin
		AssumePrime = 1;
	end	else if (num==16'd40177) begin
		AssumePrime = 1;
	end	else if (num==16'd40189) begin
		AssumePrime = 1;
	end	else if (num==16'd40193) begin
		AssumePrime = 1;
	end	else if (num==16'd40213) begin
		AssumePrime = 1;
	end	else if (num==16'd40231) begin
		AssumePrime = 1;
	end	else if (num==16'd40237) begin
		AssumePrime = 1;
	end	else if (num==16'd40241) begin
		AssumePrime = 1;
	end	else if (num==16'd40253) begin
		AssumePrime = 1;
	end	else if (num==16'd40277) begin
		AssumePrime = 1;
	end	else if (num==16'd40283) begin
		AssumePrime = 1;
	end	else if (num==16'd40289) begin
		AssumePrime = 1;
	end	else if (num==16'd40343) begin
		AssumePrime = 1;
	end	else if (num==16'd40351) begin
		AssumePrime = 1;
	end	else if (num==16'd40357) begin
		AssumePrime = 1;
	end	else if (num==16'd40361) begin
		AssumePrime = 1;
	end	else if (num==16'd40387) begin
		AssumePrime = 1;
	end	else if (num==16'd40423) begin
		AssumePrime = 1;
	end	else if (num==16'd40427) begin
		AssumePrime = 1;
	end	else if (num==16'd40429) begin
		AssumePrime = 1;
	end	else if (num==16'd40433) begin
		AssumePrime = 1;
	end	else if (num==16'd40459) begin
		AssumePrime = 1;
	end	else if (num==16'd40471) begin
		AssumePrime = 1;
	end	else if (num==16'd40483) begin
		AssumePrime = 1;
	end	else if (num==16'd40487) begin
		AssumePrime = 1;
	end	else if (num==16'd40493) begin
		AssumePrime = 1;
	end	else if (num==16'd40499) begin
		AssumePrime = 1;
	end	else if (num==16'd40507) begin
		AssumePrime = 1;
	end	else if (num==16'd40519) begin
		AssumePrime = 1;
	end	else if (num==16'd40529) begin
		AssumePrime = 1;
	end	else if (num==16'd40531) begin
		AssumePrime = 1;
	end	else if (num==16'd40543) begin
		AssumePrime = 1;
	end	else if (num==16'd40559) begin
		AssumePrime = 1;
	end	else if (num==16'd40577) begin
		AssumePrime = 1;
	end	else if (num==16'd40583) begin
		AssumePrime = 1;
	end	else if (num==16'd40591) begin
		AssumePrime = 1;
	end	else if (num==16'd40597) begin
		AssumePrime = 1;
	end	else if (num==16'd40609) begin
		AssumePrime = 1;
	end	else if (num==16'd40627) begin
		AssumePrime = 1;
	end	else if (num==16'd40637) begin
		AssumePrime = 1;
	end	else if (num==16'd40639) begin
		AssumePrime = 1;
	end	else if (num==16'd40693) begin
		AssumePrime = 1;
	end	else if (num==16'd40697) begin
		AssumePrime = 1;
	end	else if (num==16'd40699) begin
		AssumePrime = 1;
	end	else if (num==16'd40709) begin
		AssumePrime = 1;
	end	else if (num==16'd40739) begin
		AssumePrime = 1;
	end	else if (num==16'd40751) begin
		AssumePrime = 1;
	end	else if (num==16'd40759) begin
		AssumePrime = 1;
	end	else if (num==16'd40763) begin
		AssumePrime = 1;
	end	else if (num==16'd40771) begin
		AssumePrime = 1;
	end	else if (num==16'd40787) begin
		AssumePrime = 1;
	end	else if (num==16'd40801) begin
		AssumePrime = 1;
	end	else if (num==16'd40813) begin
		AssumePrime = 1;
	end	else if (num==16'd40819) begin
		AssumePrime = 1;
	end	else if (num==16'd40823) begin
		AssumePrime = 1;
	end	else if (num==16'd40829) begin
		AssumePrime = 1;
	end	else if (num==16'd40841) begin
		AssumePrime = 1;
	end	else if (num==16'd40847) begin
		AssumePrime = 1;
	end	else if (num==16'd40849) begin
		AssumePrime = 1;
	end	else if (num==16'd40853) begin
		AssumePrime = 1;
	end	else if (num==16'd40867) begin
		AssumePrime = 1;
	end	else if (num==16'd40879) begin
		AssumePrime = 1;
	end	else if (num==16'd40883) begin
		AssumePrime = 1;
	end	else if (num==16'd40897) begin
		AssumePrime = 1;
	end	else if (num==16'd40903) begin
		AssumePrime = 1;
	end	else if (num==16'd40927) begin
		AssumePrime = 1;
	end	else if (num==16'd40933) begin
		AssumePrime = 1;
	end	else if (num==16'd40939) begin
		AssumePrime = 1;
	end	else if (num==16'd40949) begin
		AssumePrime = 1;
	end	else if (num==16'd40961) begin
		AssumePrime = 1;
	end	else if (num==16'd40973) begin
		AssumePrime = 1;
	end	else if (num==16'd40993) begin
		AssumePrime = 1;
	end	else if (num==16'd41011) begin
		AssumePrime = 1;
	end	else if (num==16'd41017) begin
		AssumePrime = 1;
	end	else if (num==16'd41023) begin
		AssumePrime = 1;
	end	else if (num==16'd41039) begin
		AssumePrime = 1;
	end	else if (num==16'd41047) begin
		AssumePrime = 1;
	end	else if (num==16'd41051) begin
		AssumePrime = 1;
	end	else if (num==16'd41057) begin
		AssumePrime = 1;
	end	else if (num==16'd41077) begin
		AssumePrime = 1;
	end	else if (num==16'd41081) begin
		AssumePrime = 1;
	end	else if (num==16'd41113) begin
		AssumePrime = 1;
	end	else if (num==16'd41117) begin
		AssumePrime = 1;
	end	else if (num==16'd41131) begin
		AssumePrime = 1;
	end	else if (num==16'd41141) begin
		AssumePrime = 1;
	end	else if (num==16'd41143) begin
		AssumePrime = 1;
	end	else if (num==16'd41149) begin
		AssumePrime = 1;
	end	else if (num==16'd41161) begin
		AssumePrime = 1;
	end	else if (num==16'd41177) begin
		AssumePrime = 1;
	end	else if (num==16'd41179) begin
		AssumePrime = 1;
	end	else if (num==16'd41183) begin
		AssumePrime = 1;
	end	else if (num==16'd41189) begin
		AssumePrime = 1;
	end	else if (num==16'd41201) begin
		AssumePrime = 1;
	end	else if (num==16'd41203) begin
		AssumePrime = 1;
	end	else if (num==16'd41213) begin
		AssumePrime = 1;
	end	else if (num==16'd41221) begin
		AssumePrime = 1;
	end	else if (num==16'd41227) begin
		AssumePrime = 1;
	end	else if (num==16'd41231) begin
		AssumePrime = 1;
	end	else if (num==16'd41233) begin
		AssumePrime = 1;
	end	else if (num==16'd41243) begin
		AssumePrime = 1;
	end	else if (num==16'd41257) begin
		AssumePrime = 1;
	end	else if (num==16'd41263) begin
		AssumePrime = 1;
	end	else if (num==16'd41269) begin
		AssumePrime = 1;
	end	else if (num==16'd41281) begin
		AssumePrime = 1;
	end	else if (num==16'd41299) begin
		AssumePrime = 1;
	end	else if (num==16'd41333) begin
		AssumePrime = 1;
	end	else if (num==16'd41341) begin
		AssumePrime = 1;
	end	else if (num==16'd41351) begin
		AssumePrime = 1;
	end	else if (num==16'd41357) begin
		AssumePrime = 1;
	end	else if (num==16'd41381) begin
		AssumePrime = 1;
	end	else if (num==16'd41387) begin
		AssumePrime = 1;
	end	else if (num==16'd41389) begin
		AssumePrime = 1;
	end	else if (num==16'd41399) begin
		AssumePrime = 1;
	end	else if (num==16'd41411) begin
		AssumePrime = 1;
	end	else if (num==16'd41413) begin
		AssumePrime = 1;
	end	else if (num==16'd41443) begin
		AssumePrime = 1;
	end	else if (num==16'd41453) begin
		AssumePrime = 1;
	end	else if (num==16'd41467) begin
		AssumePrime = 1;
	end	else if (num==16'd41479) begin
		AssumePrime = 1;
	end	else if (num==16'd41491) begin
		AssumePrime = 1;
	end	else if (num==16'd41507) begin
		AssumePrime = 1;
	end	else if (num==16'd41513) begin
		AssumePrime = 1;
	end	else if (num==16'd41519) begin
		AssumePrime = 1;
	end	else if (num==16'd41521) begin
		AssumePrime = 1;
	end	else if (num==16'd41539) begin
		AssumePrime = 1;
	end	else if (num==16'd41543) begin
		AssumePrime = 1;
	end	else if (num==16'd41549) begin
		AssumePrime = 1;
	end	else if (num==16'd41579) begin
		AssumePrime = 1;
	end	else if (num==16'd41593) begin
		AssumePrime = 1;
	end	else if (num==16'd41597) begin
		AssumePrime = 1;
	end	else if (num==16'd41603) begin
		AssumePrime = 1;
	end	else if (num==16'd41609) begin
		AssumePrime = 1;
	end	else if (num==16'd41611) begin
		AssumePrime = 1;
	end	else if (num==16'd41617) begin
		AssumePrime = 1;
	end	else if (num==16'd41621) begin
		AssumePrime = 1;
	end	else if (num==16'd41627) begin
		AssumePrime = 1;
	end	else if (num==16'd41641) begin
		AssumePrime = 1;
	end	else if (num==16'd41647) begin
		AssumePrime = 1;
	end	else if (num==16'd41651) begin
		AssumePrime = 1;
	end	else if (num==16'd41659) begin
		AssumePrime = 1;
	end	else if (num==16'd41669) begin
		AssumePrime = 1;
	end	else if (num==16'd41681) begin
		AssumePrime = 1;
	end	else if (num==16'd41687) begin
		AssumePrime = 1;
	end	else if (num==16'd41719) begin
		AssumePrime = 1;
	end	else if (num==16'd41729) begin
		AssumePrime = 1;
	end	else if (num==16'd41737) begin
		AssumePrime = 1;
	end	else if (num==16'd41759) begin
		AssumePrime = 1;
	end	else if (num==16'd41761) begin
		AssumePrime = 1;
	end	else if (num==16'd41771) begin
		AssumePrime = 1;
	end	else if (num==16'd41777) begin
		AssumePrime = 1;
	end	else if (num==16'd41801) begin
		AssumePrime = 1;
	end	else if (num==16'd41809) begin
		AssumePrime = 1;
	end	else if (num==16'd41813) begin
		AssumePrime = 1;
	end	else if (num==16'd41843) begin
		AssumePrime = 1;
	end	else if (num==16'd41849) begin
		AssumePrime = 1;
	end	else if (num==16'd41851) begin
		AssumePrime = 1;
	end	else if (num==16'd41863) begin
		AssumePrime = 1;
	end	else if (num==16'd41879) begin
		AssumePrime = 1;
	end	else if (num==16'd41887) begin
		AssumePrime = 1;
	end	else if (num==16'd41893) begin
		AssumePrime = 1;
	end	else if (num==16'd41897) begin
		AssumePrime = 1;
	end	else if (num==16'd41903) begin
		AssumePrime = 1;
	end	else if (num==16'd41911) begin
		AssumePrime = 1;
	end	else if (num==16'd41927) begin
		AssumePrime = 1;
	end	else if (num==16'd41941) begin
		AssumePrime = 1;
	end	else if (num==16'd41947) begin
		AssumePrime = 1;
	end	else if (num==16'd41953) begin
		AssumePrime = 1;
	end	else if (num==16'd41957) begin
		AssumePrime = 1;
	end	else if (num==16'd41959) begin
		AssumePrime = 1;
	end	else if (num==16'd41969) begin
		AssumePrime = 1;
	end	else if (num==16'd41981) begin
		AssumePrime = 1;
	end	else if (num==16'd41983) begin
		AssumePrime = 1;
	end	else if (num==16'd41999) begin
		AssumePrime = 1;
	end	else if (num==16'd42013) begin
		AssumePrime = 1;
	end	else if (num==16'd42017) begin
		AssumePrime = 1;
	end	else if (num==16'd42019) begin
		AssumePrime = 1;
	end	else if (num==16'd42023) begin
		AssumePrime = 1;
	end	else if (num==16'd42043) begin
		AssumePrime = 1;
	end	else if (num==16'd42061) begin
		AssumePrime = 1;
	end	else if (num==16'd42071) begin
		AssumePrime = 1;
	end	else if (num==16'd42073) begin
		AssumePrime = 1;
	end	else if (num==16'd42083) begin
		AssumePrime = 1;
	end	else if (num==16'd42089) begin
		AssumePrime = 1;
	end	else if (num==16'd42101) begin
		AssumePrime = 1;
	end	else if (num==16'd42131) begin
		AssumePrime = 1;
	end	else if (num==16'd42139) begin
		AssumePrime = 1;
	end	else if (num==16'd42157) begin
		AssumePrime = 1;
	end	else if (num==16'd42169) begin
		AssumePrime = 1;
	end	else if (num==16'd42179) begin
		AssumePrime = 1;
	end	else if (num==16'd42181) begin
		AssumePrime = 1;
	end	else if (num==16'd42187) begin
		AssumePrime = 1;
	end	else if (num==16'd42193) begin
		AssumePrime = 1;
	end	else if (num==16'd42197) begin
		AssumePrime = 1;
	end	else if (num==16'd42209) begin
		AssumePrime = 1;
	end	else if (num==16'd42221) begin
		AssumePrime = 1;
	end	else if (num==16'd42223) begin
		AssumePrime = 1;
	end	else if (num==16'd42227) begin
		AssumePrime = 1;
	end	else if (num==16'd42239) begin
		AssumePrime = 1;
	end	else if (num==16'd42257) begin
		AssumePrime = 1;
	end	else if (num==16'd42281) begin
		AssumePrime = 1;
	end	else if (num==16'd42283) begin
		AssumePrime = 1;
	end	else if (num==16'd42293) begin
		AssumePrime = 1;
	end	else if (num==16'd42299) begin
		AssumePrime = 1;
	end	else if (num==16'd42307) begin
		AssumePrime = 1;
	end	else if (num==16'd42323) begin
		AssumePrime = 1;
	end	else if (num==16'd42331) begin
		AssumePrime = 1;
	end	else if (num==16'd42337) begin
		AssumePrime = 1;
	end	else if (num==16'd42349) begin
		AssumePrime = 1;
	end	else if (num==16'd42359) begin
		AssumePrime = 1;
	end	else if (num==16'd42373) begin
		AssumePrime = 1;
	end	else if (num==16'd42379) begin
		AssumePrime = 1;
	end	else if (num==16'd42391) begin
		AssumePrime = 1;
	end	else if (num==16'd42397) begin
		AssumePrime = 1;
	end	else if (num==16'd42403) begin
		AssumePrime = 1;
	end	else if (num==16'd42407) begin
		AssumePrime = 1;
	end	else if (num==16'd42409) begin
		AssumePrime = 1;
	end	else if (num==16'd42433) begin
		AssumePrime = 1;
	end	else if (num==16'd42437) begin
		AssumePrime = 1;
	end	else if (num==16'd42443) begin
		AssumePrime = 1;
	end	else if (num==16'd42451) begin
		AssumePrime = 1;
	end	else if (num==16'd42457) begin
		AssumePrime = 1;
	end	else if (num==16'd42461) begin
		AssumePrime = 1;
	end	else if (num==16'd42463) begin
		AssumePrime = 1;
	end	else if (num==16'd42467) begin
		AssumePrime = 1;
	end	else if (num==16'd42473) begin
		AssumePrime = 1;
	end	else if (num==16'd42487) begin
		AssumePrime = 1;
	end	else if (num==16'd42491) begin
		AssumePrime = 1;
	end	else if (num==16'd42499) begin
		AssumePrime = 1;
	end	else if (num==16'd42509) begin
		AssumePrime = 1;
	end	else if (num==16'd42533) begin
		AssumePrime = 1;
	end	else if (num==16'd42557) begin
		AssumePrime = 1;
	end	else if (num==16'd42569) begin
		AssumePrime = 1;
	end	else if (num==16'd42571) begin
		AssumePrime = 1;
	end	else if (num==16'd42577) begin
		AssumePrime = 1;
	end	else if (num==16'd42589) begin
		AssumePrime = 1;
	end	else if (num==16'd42611) begin
		AssumePrime = 1;
	end	else if (num==16'd42641) begin
		AssumePrime = 1;
	end	else if (num==16'd42643) begin
		AssumePrime = 1;
	end	else if (num==16'd42649) begin
		AssumePrime = 1;
	end	else if (num==16'd42667) begin
		AssumePrime = 1;
	end	else if (num==16'd42677) begin
		AssumePrime = 1;
	end	else if (num==16'd42683) begin
		AssumePrime = 1;
	end	else if (num==16'd42689) begin
		AssumePrime = 1;
	end	else if (num==16'd42697) begin
		AssumePrime = 1;
	end	else if (num==16'd42701) begin
		AssumePrime = 1;
	end	else if (num==16'd42703) begin
		AssumePrime = 1;
	end	else if (num==16'd42709) begin
		AssumePrime = 1;
	end	else if (num==16'd42719) begin
		AssumePrime = 1;
	end	else if (num==16'd42727) begin
		AssumePrime = 1;
	end	else if (num==16'd42737) begin
		AssumePrime = 1;
	end	else if (num==16'd42743) begin
		AssumePrime = 1;
	end	else if (num==16'd42751) begin
		AssumePrime = 1;
	end	else if (num==16'd42767) begin
		AssumePrime = 1;
	end	else if (num==16'd42773) begin
		AssumePrime = 1;
	end	else if (num==16'd42787) begin
		AssumePrime = 1;
	end	else if (num==16'd42793) begin
		AssumePrime = 1;
	end	else if (num==16'd42797) begin
		AssumePrime = 1;
	end	else if (num==16'd42821) begin
		AssumePrime = 1;
	end	else if (num==16'd42829) begin
		AssumePrime = 1;
	end	else if (num==16'd42839) begin
		AssumePrime = 1;
	end	else if (num==16'd42841) begin
		AssumePrime = 1;
	end	else if (num==16'd42853) begin
		AssumePrime = 1;
	end	else if (num==16'd42859) begin
		AssumePrime = 1;
	end	else if (num==16'd42863) begin
		AssumePrime = 1;
	end	else if (num==16'd42899) begin
		AssumePrime = 1;
	end	else if (num==16'd42901) begin
		AssumePrime = 1;
	end	else if (num==16'd42923) begin
		AssumePrime = 1;
	end	else if (num==16'd42929) begin
		AssumePrime = 1;
	end	else if (num==16'd42937) begin
		AssumePrime = 1;
	end	else if (num==16'd42943) begin
		AssumePrime = 1;
	end	else if (num==16'd42953) begin
		AssumePrime = 1;
	end	else if (num==16'd42961) begin
		AssumePrime = 1;
	end	else if (num==16'd42967) begin
		AssumePrime = 1;
	end	else if (num==16'd42979) begin
		AssumePrime = 1;
	end	else if (num==16'd42989) begin
		AssumePrime = 1;
	end	else if (num==16'd43003) begin
		AssumePrime = 1;
	end	else if (num==16'd43013) begin
		AssumePrime = 1;
	end	else if (num==16'd43019) begin
		AssumePrime = 1;
	end	else if (num==16'd43037) begin
		AssumePrime = 1;
	end	else if (num==16'd43049) begin
		AssumePrime = 1;
	end	else if (num==16'd43051) begin
		AssumePrime = 1;
	end	else if (num==16'd43063) begin
		AssumePrime = 1;
	end	else if (num==16'd43067) begin
		AssumePrime = 1;
	end	else if (num==16'd43093) begin
		AssumePrime = 1;
	end	else if (num==16'd43103) begin
		AssumePrime = 1;
	end	else if (num==16'd43117) begin
		AssumePrime = 1;
	end	else if (num==16'd43133) begin
		AssumePrime = 1;
	end	else if (num==16'd43151) begin
		AssumePrime = 1;
	end	else if (num==16'd43159) begin
		AssumePrime = 1;
	end	else if (num==16'd43177) begin
		AssumePrime = 1;
	end	else if (num==16'd43189) begin
		AssumePrime = 1;
	end	else if (num==16'd43201) begin
		AssumePrime = 1;
	end	else if (num==16'd43207) begin
		AssumePrime = 1;
	end	else if (num==16'd43223) begin
		AssumePrime = 1;
	end	else if (num==16'd43237) begin
		AssumePrime = 1;
	end	else if (num==16'd43261) begin
		AssumePrime = 1;
	end	else if (num==16'd43271) begin
		AssumePrime = 1;
	end	else if (num==16'd43283) begin
		AssumePrime = 1;
	end	else if (num==16'd43291) begin
		AssumePrime = 1;
	end	else if (num==16'd43313) begin
		AssumePrime = 1;
	end	else if (num==16'd43319) begin
		AssumePrime = 1;
	end	else if (num==16'd43321) begin
		AssumePrime = 1;
	end	else if (num==16'd43331) begin
		AssumePrime = 1;
	end	else if (num==16'd43391) begin
		AssumePrime = 1;
	end	else if (num==16'd43397) begin
		AssumePrime = 1;
	end	else if (num==16'd43399) begin
		AssumePrime = 1;
	end	else if (num==16'd43403) begin
		AssumePrime = 1;
	end	else if (num==16'd43411) begin
		AssumePrime = 1;
	end	else if (num==16'd43427) begin
		AssumePrime = 1;
	end	else if (num==16'd43441) begin
		AssumePrime = 1;
	end	else if (num==16'd43451) begin
		AssumePrime = 1;
	end	else if (num==16'd43457) begin
		AssumePrime = 1;
	end	else if (num==16'd43481) begin
		AssumePrime = 1;
	end	else if (num==16'd43487) begin
		AssumePrime = 1;
	end	else if (num==16'd43499) begin
		AssumePrime = 1;
	end	else if (num==16'd43517) begin
		AssumePrime = 1;
	end	else if (num==16'd43541) begin
		AssumePrime = 1;
	end	else if (num==16'd43543) begin
		AssumePrime = 1;
	end	else if (num==16'd43573) begin
		AssumePrime = 1;
	end	else if (num==16'd43577) begin
		AssumePrime = 1;
	end	else if (num==16'd43579) begin
		AssumePrime = 1;
	end	else if (num==16'd43591) begin
		AssumePrime = 1;
	end	else if (num==16'd43597) begin
		AssumePrime = 1;
	end	else if (num==16'd43607) begin
		AssumePrime = 1;
	end	else if (num==16'd43609) begin
		AssumePrime = 1;
	end	else if (num==16'd43613) begin
		AssumePrime = 1;
	end	else if (num==16'd43627) begin
		AssumePrime = 1;
	end	else if (num==16'd43633) begin
		AssumePrime = 1;
	end	else if (num==16'd43649) begin
		AssumePrime = 1;
	end	else if (num==16'd43651) begin
		AssumePrime = 1;
	end	else if (num==16'd43661) begin
		AssumePrime = 1;
	end	else if (num==16'd43669) begin
		AssumePrime = 1;
	end	else if (num==16'd43691) begin
		AssumePrime = 1;
	end	else if (num==16'd43711) begin
		AssumePrime = 1;
	end	else if (num==16'd43717) begin
		AssumePrime = 1;
	end	else if (num==16'd43721) begin
		AssumePrime = 1;
	end	else if (num==16'd43753) begin
		AssumePrime = 1;
	end	else if (num==16'd43759) begin
		AssumePrime = 1;
	end	else if (num==16'd43777) begin
		AssumePrime = 1;
	end	else if (num==16'd43781) begin
		AssumePrime = 1;
	end	else if (num==16'd43783) begin
		AssumePrime = 1;
	end	else if (num==16'd43787) begin
		AssumePrime = 1;
	end	else if (num==16'd43789) begin
		AssumePrime = 1;
	end	else if (num==16'd43793) begin
		AssumePrime = 1;
	end	else if (num==16'd43801) begin
		AssumePrime = 1;
	end	else if (num==16'd43853) begin
		AssumePrime = 1;
	end	else if (num==16'd43867) begin
		AssumePrime = 1;
	end	else if (num==16'd43889) begin
		AssumePrime = 1;
	end	else if (num==16'd43891) begin
		AssumePrime = 1;
	end	else if (num==16'd43913) begin
		AssumePrime = 1;
	end	else if (num==16'd43933) begin
		AssumePrime = 1;
	end	else if (num==16'd43943) begin
		AssumePrime = 1;
	end	else if (num==16'd43951) begin
		AssumePrime = 1;
	end	else if (num==16'd43961) begin
		AssumePrime = 1;
	end	else if (num==16'd43963) begin
		AssumePrime = 1;
	end	else if (num==16'd43969) begin
		AssumePrime = 1;
	end	else if (num==16'd43973) begin
		AssumePrime = 1;
	end	else if (num==16'd43987) begin
		AssumePrime = 1;
	end	else if (num==16'd43991) begin
		AssumePrime = 1;
	end	else if (num==16'd43997) begin
		AssumePrime = 1;
	end	else if (num==16'd44017) begin
		AssumePrime = 1;
	end	else if (num==16'd44021) begin
		AssumePrime = 1;
	end	else if (num==16'd44027) begin
		AssumePrime = 1;
	end	else if (num==16'd44029) begin
		AssumePrime = 1;
	end	else if (num==16'd44041) begin
		AssumePrime = 1;
	end	else if (num==16'd44053) begin
		AssumePrime = 1;
	end	else if (num==16'd44059) begin
		AssumePrime = 1;
	end	else if (num==16'd44071) begin
		AssumePrime = 1;
	end	else if (num==16'd44087) begin
		AssumePrime = 1;
	end	else if (num==16'd44089) begin
		AssumePrime = 1;
	end	else if (num==16'd44101) begin
		AssumePrime = 1;
	end	else if (num==16'd44111) begin
		AssumePrime = 1;
	end	else if (num==16'd44119) begin
		AssumePrime = 1;
	end	else if (num==16'd44123) begin
		AssumePrime = 1;
	end	else if (num==16'd44129) begin
		AssumePrime = 1;
	end	else if (num==16'd44131) begin
		AssumePrime = 1;
	end	else if (num==16'd44159) begin
		AssumePrime = 1;
	end	else if (num==16'd44171) begin
		AssumePrime = 1;
	end	else if (num==16'd44179) begin
		AssumePrime = 1;
	end	else if (num==16'd44189) begin
		AssumePrime = 1;
	end	else if (num==16'd44201) begin
		AssumePrime = 1;
	end	else if (num==16'd44203) begin
		AssumePrime = 1;
	end	else if (num==16'd44207) begin
		AssumePrime = 1;
	end	else if (num==16'd44221) begin
		AssumePrime = 1;
	end	else if (num==16'd44249) begin
		AssumePrime = 1;
	end	else if (num==16'd44257) begin
		AssumePrime = 1;
	end	else if (num==16'd44263) begin
		AssumePrime = 1;
	end	else if (num==16'd44267) begin
		AssumePrime = 1;
	end	else if (num==16'd44269) begin
		AssumePrime = 1;
	end	else if (num==16'd44273) begin
		AssumePrime = 1;
	end	else if (num==16'd44279) begin
		AssumePrime = 1;
	end	else if (num==16'd44281) begin
		AssumePrime = 1;
	end	else if (num==16'd44293) begin
		AssumePrime = 1;
	end	else if (num==16'd44351) begin
		AssumePrime = 1;
	end	else if (num==16'd44357) begin
		AssumePrime = 1;
	end	else if (num==16'd44371) begin
		AssumePrime = 1;
	end	else if (num==16'd44381) begin
		AssumePrime = 1;
	end	else if (num==16'd44383) begin
		AssumePrime = 1;
	end	else if (num==16'd44389) begin
		AssumePrime = 1;
	end	else if (num==16'd44417) begin
		AssumePrime = 1;
	end	else if (num==16'd44449) begin
		AssumePrime = 1;
	end	else if (num==16'd44453) begin
		AssumePrime = 1;
	end	else if (num==16'd44483) begin
		AssumePrime = 1;
	end	else if (num==16'd44491) begin
		AssumePrime = 1;
	end	else if (num==16'd44497) begin
		AssumePrime = 1;
	end	else if (num==16'd44501) begin
		AssumePrime = 1;
	end	else if (num==16'd44507) begin
		AssumePrime = 1;
	end	else if (num==16'd44519) begin
		AssumePrime = 1;
	end	else if (num==16'd44531) begin
		AssumePrime = 1;
	end	else if (num==16'd44533) begin
		AssumePrime = 1;
	end	else if (num==16'd44537) begin
		AssumePrime = 1;
	end	else if (num==16'd44543) begin
		AssumePrime = 1;
	end	else if (num==16'd44549) begin
		AssumePrime = 1;
	end	else if (num==16'd44563) begin
		AssumePrime = 1;
	end	else if (num==16'd44579) begin
		AssumePrime = 1;
	end	else if (num==16'd44587) begin
		AssumePrime = 1;
	end	else if (num==16'd44617) begin
		AssumePrime = 1;
	end	else if (num==16'd44621) begin
		AssumePrime = 1;
	end	else if (num==16'd44623) begin
		AssumePrime = 1;
	end	else if (num==16'd44633) begin
		AssumePrime = 1;
	end	else if (num==16'd44641) begin
		AssumePrime = 1;
	end	else if (num==16'd44647) begin
		AssumePrime = 1;
	end	else if (num==16'd44651) begin
		AssumePrime = 1;
	end	else if (num==16'd44657) begin
		AssumePrime = 1;
	end	else if (num==16'd44683) begin
		AssumePrime = 1;
	end	else if (num==16'd44687) begin
		AssumePrime = 1;
	end	else if (num==16'd44699) begin
		AssumePrime = 1;
	end	else if (num==16'd44701) begin
		AssumePrime = 1;
	end	else if (num==16'd44711) begin
		AssumePrime = 1;
	end	else if (num==16'd44729) begin
		AssumePrime = 1;
	end	else if (num==16'd44741) begin
		AssumePrime = 1;
	end	else if (num==16'd44753) begin
		AssumePrime = 1;
	end	else if (num==16'd44771) begin
		AssumePrime = 1;
	end	else if (num==16'd44773) begin
		AssumePrime = 1;
	end	else if (num==16'd44777) begin
		AssumePrime = 1;
	end	else if (num==16'd44789) begin
		AssumePrime = 1;
	end	else if (num==16'd44797) begin
		AssumePrime = 1;
	end	else if (num==16'd44809) begin
		AssumePrime = 1;
	end	else if (num==16'd44819) begin
		AssumePrime = 1;
	end	else if (num==16'd44839) begin
		AssumePrime = 1;
	end	else if (num==16'd44843) begin
		AssumePrime = 1;
	end	else if (num==16'd44851) begin
		AssumePrime = 1;
	end	else if (num==16'd44867) begin
		AssumePrime = 1;
	end	else if (num==16'd44879) begin
		AssumePrime = 1;
	end	else if (num==16'd44887) begin
		AssumePrime = 1;
	end	else if (num==16'd44893) begin
		AssumePrime = 1;
	end	else if (num==16'd44909) begin
		AssumePrime = 1;
	end	else if (num==16'd44917) begin
		AssumePrime = 1;
	end	else if (num==16'd44927) begin
		AssumePrime = 1;
	end	else if (num==16'd44939) begin
		AssumePrime = 1;
	end	else if (num==16'd44953) begin
		AssumePrime = 1;
	end	else if (num==16'd44959) begin
		AssumePrime = 1;
	end	else if (num==16'd44963) begin
		AssumePrime = 1;
	end	else if (num==16'd44971) begin
		AssumePrime = 1;
	end	else if (num==16'd44983) begin
		AssumePrime = 1;
	end	else if (num==16'd44987) begin
		AssumePrime = 1;
	end	else if (num==16'd45007) begin
		AssumePrime = 1;
	end	else if (num==16'd45013) begin
		AssumePrime = 1;
	end	else if (num==16'd45053) begin
		AssumePrime = 1;
	end	else if (num==16'd45061) begin
		AssumePrime = 1;
	end	else if (num==16'd45077) begin
		AssumePrime = 1;
	end	else if (num==16'd45083) begin
		AssumePrime = 1;
	end	else if (num==16'd45119) begin
		AssumePrime = 1;
	end	else if (num==16'd45121) begin
		AssumePrime = 1;
	end	else if (num==16'd45127) begin
		AssumePrime = 1;
	end	else if (num==16'd45131) begin
		AssumePrime = 1;
	end	else if (num==16'd45137) begin
		AssumePrime = 1;
	end	else if (num==16'd45139) begin
		AssumePrime = 1;
	end	else if (num==16'd45161) begin
		AssumePrime = 1;
	end	else if (num==16'd45179) begin
		AssumePrime = 1;
	end	else if (num==16'd45181) begin
		AssumePrime = 1;
	end	else if (num==16'd45191) begin
		AssumePrime = 1;
	end	else if (num==16'd45197) begin
		AssumePrime = 1;
	end	else if (num==16'd45233) begin
		AssumePrime = 1;
	end	else if (num==16'd45247) begin
		AssumePrime = 1;
	end	else if (num==16'd45259) begin
		AssumePrime = 1;
	end	else if (num==16'd45263) begin
		AssumePrime = 1;
	end	else if (num==16'd45281) begin
		AssumePrime = 1;
	end	else if (num==16'd45289) begin
		AssumePrime = 1;
	end	else if (num==16'd45293) begin
		AssumePrime = 1;
	end	else if (num==16'd45307) begin
		AssumePrime = 1;
	end	else if (num==16'd45317) begin
		AssumePrime = 1;
	end	else if (num==16'd45319) begin
		AssumePrime = 1;
	end	else if (num==16'd45329) begin
		AssumePrime = 1;
	end	else if (num==16'd45337) begin
		AssumePrime = 1;
	end	else if (num==16'd45341) begin
		AssumePrime = 1;
	end	else if (num==16'd45343) begin
		AssumePrime = 1;
	end	else if (num==16'd45361) begin
		AssumePrime = 1;
	end	else if (num==16'd45377) begin
		AssumePrime = 1;
	end	else if (num==16'd45389) begin
		AssumePrime = 1;
	end	else if (num==16'd45403) begin
		AssumePrime = 1;
	end	else if (num==16'd45413) begin
		AssumePrime = 1;
	end	else if (num==16'd45427) begin
		AssumePrime = 1;
	end	else if (num==16'd45433) begin
		AssumePrime = 1;
	end	else if (num==16'd45439) begin
		AssumePrime = 1;
	end	else if (num==16'd45481) begin
		AssumePrime = 1;
	end	else if (num==16'd45491) begin
		AssumePrime = 1;
	end	else if (num==16'd45497) begin
		AssumePrime = 1;
	end	else if (num==16'd45503) begin
		AssumePrime = 1;
	end	else if (num==16'd45523) begin
		AssumePrime = 1;
	end	else if (num==16'd45533) begin
		AssumePrime = 1;
	end	else if (num==16'd45541) begin
		AssumePrime = 1;
	end	else if (num==16'd45553) begin
		AssumePrime = 1;
	end	else if (num==16'd45557) begin
		AssumePrime = 1;
	end	else if (num==16'd45569) begin
		AssumePrime = 1;
	end	else if (num==16'd45587) begin
		AssumePrime = 1;
	end	else if (num==16'd45589) begin
		AssumePrime = 1;
	end	else if (num==16'd45599) begin
		AssumePrime = 1;
	end	else if (num==16'd45613) begin
		AssumePrime = 1;
	end	else if (num==16'd45631) begin
		AssumePrime = 1;
	end	else if (num==16'd45641) begin
		AssumePrime = 1;
	end	else if (num==16'd45659) begin
		AssumePrime = 1;
	end	else if (num==16'd45667) begin
		AssumePrime = 1;
	end	else if (num==16'd45673) begin
		AssumePrime = 1;
	end	else if (num==16'd45677) begin
		AssumePrime = 1;
	end	else if (num==16'd45691) begin
		AssumePrime = 1;
	end	else if (num==16'd45697) begin
		AssumePrime = 1;
	end	else if (num==16'd45707) begin
		AssumePrime = 1;
	end	else if (num==16'd45737) begin
		AssumePrime = 1;
	end	else if (num==16'd45751) begin
		AssumePrime = 1;
	end	else if (num==16'd45757) begin
		AssumePrime = 1;
	end	else if (num==16'd45763) begin
		AssumePrime = 1;
	end	else if (num==16'd45767) begin
		AssumePrime = 1;
	end	else if (num==16'd45779) begin
		AssumePrime = 1;
	end	else if (num==16'd45817) begin
		AssumePrime = 1;
	end	else if (num==16'd45821) begin
		AssumePrime = 1;
	end	else if (num==16'd45823) begin
		AssumePrime = 1;
	end	else if (num==16'd45827) begin
		AssumePrime = 1;
	end	else if (num==16'd45833) begin
		AssumePrime = 1;
	end	else if (num==16'd45841) begin
		AssumePrime = 1;
	end	else if (num==16'd45853) begin
		AssumePrime = 1;
	end	else if (num==16'd45863) begin
		AssumePrime = 1;
	end	else if (num==16'd45869) begin
		AssumePrime = 1;
	end	else if (num==16'd45887) begin
		AssumePrime = 1;
	end	else if (num==16'd45893) begin
		AssumePrime = 1;
	end	else if (num==16'd45943) begin
		AssumePrime = 1;
	end	else if (num==16'd45949) begin
		AssumePrime = 1;
	end	else if (num==16'd45953) begin
		AssumePrime = 1;
	end	else if (num==16'd45959) begin
		AssumePrime = 1;
	end	else if (num==16'd45971) begin
		AssumePrime = 1;
	end	else if (num==16'd45979) begin
		AssumePrime = 1;
	end	else if (num==16'd45989) begin
		AssumePrime = 1;
	end	else if (num==16'd46021) begin
		AssumePrime = 1;
	end	else if (num==16'd46027) begin
		AssumePrime = 1;
	end	else if (num==16'd46049) begin
		AssumePrime = 1;
	end	else if (num==16'd46051) begin
		AssumePrime = 1;
	end	else if (num==16'd46061) begin
		AssumePrime = 1;
	end	else if (num==16'd46073) begin
		AssumePrime = 1;
	end	else if (num==16'd46091) begin
		AssumePrime = 1;
	end	else if (num==16'd46093) begin
		AssumePrime = 1;
	end	else if (num==16'd46099) begin
		AssumePrime = 1;
	end	else if (num==16'd46103) begin
		AssumePrime = 1;
	end	else if (num==16'd46133) begin
		AssumePrime = 1;
	end	else if (num==16'd46141) begin
		AssumePrime = 1;
	end	else if (num==16'd46147) begin
		AssumePrime = 1;
	end	else if (num==16'd46153) begin
		AssumePrime = 1;
	end	else if (num==16'd46171) begin
		AssumePrime = 1;
	end	else if (num==16'd46181) begin
		AssumePrime = 1;
	end	else if (num==16'd46183) begin
		AssumePrime = 1;
	end	else if (num==16'd46187) begin
		AssumePrime = 1;
	end	else if (num==16'd46199) begin
		AssumePrime = 1;
	end	else if (num==16'd46219) begin
		AssumePrime = 1;
	end	else if (num==16'd46229) begin
		AssumePrime = 1;
	end	else if (num==16'd46237) begin
		AssumePrime = 1;
	end	else if (num==16'd46261) begin
		AssumePrime = 1;
	end	else if (num==16'd46271) begin
		AssumePrime = 1;
	end	else if (num==16'd46273) begin
		AssumePrime = 1;
	end	else if (num==16'd46279) begin
		AssumePrime = 1;
	end	else if (num==16'd46301) begin
		AssumePrime = 1;
	end	else if (num==16'd46307) begin
		AssumePrime = 1;
	end	else if (num==16'd46309) begin
		AssumePrime = 1;
	end	else if (num==16'd46327) begin
		AssumePrime = 1;
	end	else if (num==16'd46337) begin
		AssumePrime = 1;
	end	else if (num==16'd46349) begin
		AssumePrime = 1;
	end	else if (num==16'd46351) begin
		AssumePrime = 1;
	end	else if (num==16'd46381) begin
		AssumePrime = 1;
	end	else if (num==16'd46399) begin
		AssumePrime = 1;
	end	else if (num==16'd46411) begin
		AssumePrime = 1;
	end	else if (num==16'd46439) begin
		AssumePrime = 1;
	end	else if (num==16'd46441) begin
		AssumePrime = 1;
	end	else if (num==16'd46447) begin
		AssumePrime = 1;
	end	else if (num==16'd46451) begin
		AssumePrime = 1;
	end	else if (num==16'd46457) begin
		AssumePrime = 1;
	end	else if (num==16'd46471) begin
		AssumePrime = 1;
	end	else if (num==16'd46477) begin
		AssumePrime = 1;
	end	else if (num==16'd46489) begin
		AssumePrime = 1;
	end	else if (num==16'd46499) begin
		AssumePrime = 1;
	end	else if (num==16'd46507) begin
		AssumePrime = 1;
	end	else if (num==16'd46511) begin
		AssumePrime = 1;
	end	else if (num==16'd46523) begin
		AssumePrime = 1;
	end	else if (num==16'd46549) begin
		AssumePrime = 1;
	end	else if (num==16'd46559) begin
		AssumePrime = 1;
	end	else if (num==16'd46567) begin
		AssumePrime = 1;
	end	else if (num==16'd46573) begin
		AssumePrime = 1;
	end	else if (num==16'd46589) begin
		AssumePrime = 1;
	end	else if (num==16'd46591) begin
		AssumePrime = 1;
	end	else if (num==16'd46601) begin
		AssumePrime = 1;
	end	else if (num==16'd46619) begin
		AssumePrime = 1;
	end	else if (num==16'd46633) begin
		AssumePrime = 1;
	end	else if (num==16'd46639) begin
		AssumePrime = 1;
	end	else if (num==16'd46643) begin
		AssumePrime = 1;
	end	else if (num==16'd46649) begin
		AssumePrime = 1;
	end	else if (num==16'd46663) begin
		AssumePrime = 1;
	end	else if (num==16'd46679) begin
		AssumePrime = 1;
	end	else if (num==16'd46681) begin
		AssumePrime = 1;
	end	else if (num==16'd46687) begin
		AssumePrime = 1;
	end	else if (num==16'd46691) begin
		AssumePrime = 1;
	end	else if (num==16'd46703) begin
		AssumePrime = 1;
	end	else if (num==16'd46723) begin
		AssumePrime = 1;
	end	else if (num==16'd46727) begin
		AssumePrime = 1;
	end	else if (num==16'd46747) begin
		AssumePrime = 1;
	end	else if (num==16'd46751) begin
		AssumePrime = 1;
	end	else if (num==16'd46757) begin
		AssumePrime = 1;
	end	else if (num==16'd46769) begin
		AssumePrime = 1;
	end	else if (num==16'd46771) begin
		AssumePrime = 1;
	end	else if (num==16'd46807) begin
		AssumePrime = 1;
	end	else if (num==16'd46811) begin
		AssumePrime = 1;
	end	else if (num==16'd46817) begin
		AssumePrime = 1;
	end	else if (num==16'd46819) begin
		AssumePrime = 1;
	end	else if (num==16'd46829) begin
		AssumePrime = 1;
	end	else if (num==16'd46831) begin
		AssumePrime = 1;
	end	else if (num==16'd46853) begin
		AssumePrime = 1;
	end	else if (num==16'd46861) begin
		AssumePrime = 1;
	end	else if (num==16'd46867) begin
		AssumePrime = 1;
	end	else if (num==16'd46877) begin
		AssumePrime = 1;
	end	else if (num==16'd46889) begin
		AssumePrime = 1;
	end	else if (num==16'd46901) begin
		AssumePrime = 1;
	end	else if (num==16'd46919) begin
		AssumePrime = 1;
	end	else if (num==16'd46933) begin
		AssumePrime = 1;
	end	else if (num==16'd46957) begin
		AssumePrime = 1;
	end	else if (num==16'd46993) begin
		AssumePrime = 1;
	end	else if (num==16'd46997) begin
		AssumePrime = 1;
	end	else if (num==16'd47017) begin
		AssumePrime = 1;
	end	else if (num==16'd47041) begin
		AssumePrime = 1;
	end	else if (num==16'd47051) begin
		AssumePrime = 1;
	end	else if (num==16'd47057) begin
		AssumePrime = 1;
	end	else if (num==16'd47059) begin
		AssumePrime = 1;
	end	else if (num==16'd47087) begin
		AssumePrime = 1;
	end	else if (num==16'd47093) begin
		AssumePrime = 1;
	end	else if (num==16'd47111) begin
		AssumePrime = 1;
	end	else if (num==16'd47119) begin
		AssumePrime = 1;
	end	else if (num==16'd47123) begin
		AssumePrime = 1;
	end	else if (num==16'd47129) begin
		AssumePrime = 1;
	end	else if (num==16'd47137) begin
		AssumePrime = 1;
	end	else if (num==16'd47143) begin
		AssumePrime = 1;
	end	else if (num==16'd47147) begin
		AssumePrime = 1;
	end	else if (num==16'd47149) begin
		AssumePrime = 1;
	end	else if (num==16'd47161) begin
		AssumePrime = 1;
	end	else if (num==16'd47189) begin
		AssumePrime = 1;
	end	else if (num==16'd47207) begin
		AssumePrime = 1;
	end	else if (num==16'd47221) begin
		AssumePrime = 1;
	end	else if (num==16'd47237) begin
		AssumePrime = 1;
	end	else if (num==16'd47251) begin
		AssumePrime = 1;
	end	else if (num==16'd47269) begin
		AssumePrime = 1;
	end	else if (num==16'd47279) begin
		AssumePrime = 1;
	end	else if (num==16'd47287) begin
		AssumePrime = 1;
	end	else if (num==16'd47293) begin
		AssumePrime = 1;
	end	else if (num==16'd47297) begin
		AssumePrime = 1;
	end	else if (num==16'd47303) begin
		AssumePrime = 1;
	end	else if (num==16'd47309) begin
		AssumePrime = 1;
	end	else if (num==16'd47317) begin
		AssumePrime = 1;
	end	else if (num==16'd47339) begin
		AssumePrime = 1;
	end	else if (num==16'd47351) begin
		AssumePrime = 1;
	end	else if (num==16'd47353) begin
		AssumePrime = 1;
	end	else if (num==16'd47363) begin
		AssumePrime = 1;
	end	else if (num==16'd47381) begin
		AssumePrime = 1;
	end	else if (num==16'd47387) begin
		AssumePrime = 1;
	end	else if (num==16'd47389) begin
		AssumePrime = 1;
	end	else if (num==16'd47407) begin
		AssumePrime = 1;
	end	else if (num==16'd47417) begin
		AssumePrime = 1;
	end	else if (num==16'd47419) begin
		AssumePrime = 1;
	end	else if (num==16'd47431) begin
		AssumePrime = 1;
	end	else if (num==16'd47441) begin
		AssumePrime = 1;
	end	else if (num==16'd47459) begin
		AssumePrime = 1;
	end	else if (num==16'd47491) begin
		AssumePrime = 1;
	end	else if (num==16'd47497) begin
		AssumePrime = 1;
	end	else if (num==16'd47501) begin
		AssumePrime = 1;
	end	else if (num==16'd47507) begin
		AssumePrime = 1;
	end	else if (num==16'd47513) begin
		AssumePrime = 1;
	end	else if (num==16'd47521) begin
		AssumePrime = 1;
	end	else if (num==16'd47527) begin
		AssumePrime = 1;
	end	else if (num==16'd47533) begin
		AssumePrime = 1;
	end	else if (num==16'd47543) begin
		AssumePrime = 1;
	end	else if (num==16'd47563) begin
		AssumePrime = 1;
	end	else if (num==16'd47569) begin
		AssumePrime = 1;
	end	else if (num==16'd47581) begin
		AssumePrime = 1;
	end	else if (num==16'd47591) begin
		AssumePrime = 1;
	end	else if (num==16'd47599) begin
		AssumePrime = 1;
	end	else if (num==16'd47609) begin
		AssumePrime = 1;
	end	else if (num==16'd47623) begin
		AssumePrime = 1;
	end	else if (num==16'd47629) begin
		AssumePrime = 1;
	end	else if (num==16'd47639) begin
		AssumePrime = 1;
	end	else if (num==16'd47653) begin
		AssumePrime = 1;
	end	else if (num==16'd47657) begin
		AssumePrime = 1;
	end	else if (num==16'd47659) begin
		AssumePrime = 1;
	end	else if (num==16'd47681) begin
		AssumePrime = 1;
	end	else if (num==16'd47699) begin
		AssumePrime = 1;
	end	else if (num==16'd47701) begin
		AssumePrime = 1;
	end	else if (num==16'd47711) begin
		AssumePrime = 1;
	end	else if (num==16'd47713) begin
		AssumePrime = 1;
	end	else if (num==16'd47717) begin
		AssumePrime = 1;
	end	else if (num==16'd47737) begin
		AssumePrime = 1;
	end	else if (num==16'd47741) begin
		AssumePrime = 1;
	end	else if (num==16'd47743) begin
		AssumePrime = 1;
	end	else if (num==16'd47777) begin
		AssumePrime = 1;
	end	else if (num==16'd47779) begin
		AssumePrime = 1;
	end	else if (num==16'd47791) begin
		AssumePrime = 1;
	end	else if (num==16'd47797) begin
		AssumePrime = 1;
	end	else if (num==16'd47807) begin
		AssumePrime = 1;
	end	else if (num==16'd47809) begin
		AssumePrime = 1;
	end	else if (num==16'd47819) begin
		AssumePrime = 1;
	end	else if (num==16'd47837) begin
		AssumePrime = 1;
	end	else if (num==16'd47843) begin
		AssumePrime = 1;
	end	else if (num==16'd47857) begin
		AssumePrime = 1;
	end	else if (num==16'd47869) begin
		AssumePrime = 1;
	end	else if (num==16'd47881) begin
		AssumePrime = 1;
	end	else if (num==16'd47903) begin
		AssumePrime = 1;
	end	else if (num==16'd47911) begin
		AssumePrime = 1;
	end	else if (num==16'd47917) begin
		AssumePrime = 1;
	end	else if (num==16'd47933) begin
		AssumePrime = 1;
	end	else if (num==16'd47939) begin
		AssumePrime = 1;
	end	else if (num==16'd47947) begin
		AssumePrime = 1;
	end	else if (num==16'd47951) begin
		AssumePrime = 1;
	end	else if (num==16'd47963) begin
		AssumePrime = 1;
	end	else if (num==16'd47969) begin
		AssumePrime = 1;
	end	else if (num==16'd47977) begin
		AssumePrime = 1;
	end	else if (num==16'd47981) begin
		AssumePrime = 1;
	end	else if (num==16'd48017) begin
		AssumePrime = 1;
	end	else if (num==16'd48023) begin
		AssumePrime = 1;
	end	else if (num==16'd48029) begin
		AssumePrime = 1;
	end	else if (num==16'd48049) begin
		AssumePrime = 1;
	end	else if (num==16'd48073) begin
		AssumePrime = 1;
	end	else if (num==16'd48079) begin
		AssumePrime = 1;
	end	else if (num==16'd48091) begin
		AssumePrime = 1;
	end	else if (num==16'd48109) begin
		AssumePrime = 1;
	end	else if (num==16'd48119) begin
		AssumePrime = 1;
	end	else if (num==16'd48121) begin
		AssumePrime = 1;
	end	else if (num==16'd48131) begin
		AssumePrime = 1;
	end	else if (num==16'd48157) begin
		AssumePrime = 1;
	end	else if (num==16'd48163) begin
		AssumePrime = 1;
	end	else if (num==16'd48179) begin
		AssumePrime = 1;
	end	else if (num==16'd48187) begin
		AssumePrime = 1;
	end	else if (num==16'd48193) begin
		AssumePrime = 1;
	end	else if (num==16'd48197) begin
		AssumePrime = 1;
	end	else if (num==16'd48221) begin
		AssumePrime = 1;
	end	else if (num==16'd48239) begin
		AssumePrime = 1;
	end	else if (num==16'd48247) begin
		AssumePrime = 1;
	end	else if (num==16'd48259) begin
		AssumePrime = 1;
	end	else if (num==16'd48271) begin
		AssumePrime = 1;
	end	else if (num==16'd48281) begin
		AssumePrime = 1;
	end	else if (num==16'd48299) begin
		AssumePrime = 1;
	end	else if (num==16'd48311) begin
		AssumePrime = 1;
	end	else if (num==16'd48313) begin
		AssumePrime = 1;
	end	else if (num==16'd48337) begin
		AssumePrime = 1;
	end	else if (num==16'd48341) begin
		AssumePrime = 1;
	end	else if (num==16'd48353) begin
		AssumePrime = 1;
	end	else if (num==16'd48371) begin
		AssumePrime = 1;
	end	else if (num==16'd48383) begin
		AssumePrime = 1;
	end	else if (num==16'd48397) begin
		AssumePrime = 1;
	end	else if (num==16'd48407) begin
		AssumePrime = 1;
	end	else if (num==16'd48409) begin
		AssumePrime = 1;
	end	else if (num==16'd48413) begin
		AssumePrime = 1;
	end	else if (num==16'd48437) begin
		AssumePrime = 1;
	end	else if (num==16'd48449) begin
		AssumePrime = 1;
	end	else if (num==16'd48463) begin
		AssumePrime = 1;
	end	else if (num==16'd48473) begin
		AssumePrime = 1;
	end	else if (num==16'd48479) begin
		AssumePrime = 1;
	end	else if (num==16'd48481) begin
		AssumePrime = 1;
	end	else if (num==16'd48487) begin
		AssumePrime = 1;
	end	else if (num==16'd48491) begin
		AssumePrime = 1;
	end	else if (num==16'd48497) begin
		AssumePrime = 1;
	end	else if (num==16'd48523) begin
		AssumePrime = 1;
	end	else if (num==16'd48527) begin
		AssumePrime = 1;
	end	else if (num==16'd48533) begin
		AssumePrime = 1;
	end	else if (num==16'd48539) begin
		AssumePrime = 1;
	end	else if (num==16'd48541) begin
		AssumePrime = 1;
	end	else if (num==16'd48563) begin
		AssumePrime = 1;
	end	else if (num==16'd48571) begin
		AssumePrime = 1;
	end	else if (num==16'd48589) begin
		AssumePrime = 1;
	end	else if (num==16'd48593) begin
		AssumePrime = 1;
	end	else if (num==16'd48611) begin
		AssumePrime = 1;
	end	else if (num==16'd48619) begin
		AssumePrime = 1;
	end	else if (num==16'd48623) begin
		AssumePrime = 1;
	end	else if (num==16'd48647) begin
		AssumePrime = 1;
	end	else if (num==16'd48649) begin
		AssumePrime = 1;
	end	else if (num==16'd48661) begin
		AssumePrime = 1;
	end	else if (num==16'd48673) begin
		AssumePrime = 1;
	end	else if (num==16'd48677) begin
		AssumePrime = 1;
	end	else if (num==16'd48679) begin
		AssumePrime = 1;
	end	else if (num==16'd48731) begin
		AssumePrime = 1;
	end	else if (num==16'd48733) begin
		AssumePrime = 1;
	end	else if (num==16'd48751) begin
		AssumePrime = 1;
	end	else if (num==16'd48757) begin
		AssumePrime = 1;
	end	else if (num==16'd48761) begin
		AssumePrime = 1;
	end	else if (num==16'd48767) begin
		AssumePrime = 1;
	end	else if (num==16'd48779) begin
		AssumePrime = 1;
	end	else if (num==16'd48781) begin
		AssumePrime = 1;
	end	else if (num==16'd48787) begin
		AssumePrime = 1;
	end	else if (num==16'd48799) begin
		AssumePrime = 1;
	end	else if (num==16'd48809) begin
		AssumePrime = 1;
	end	else if (num==16'd48817) begin
		AssumePrime = 1;
	end	else if (num==16'd48821) begin
		AssumePrime = 1;
	end	else if (num==16'd48823) begin
		AssumePrime = 1;
	end	else if (num==16'd48847) begin
		AssumePrime = 1;
	end	else if (num==16'd48857) begin
		AssumePrime = 1;
	end	else if (num==16'd48859) begin
		AssumePrime = 1;
	end	else if (num==16'd48869) begin
		AssumePrime = 1;
	end	else if (num==16'd48871) begin
		AssumePrime = 1;
	end	else if (num==16'd48883) begin
		AssumePrime = 1;
	end	else if (num==16'd48889) begin
		AssumePrime = 1;
	end	else if (num==16'd48907) begin
		AssumePrime = 1;
	end	else if (num==16'd48947) begin
		AssumePrime = 1;
	end	else if (num==16'd48953) begin
		AssumePrime = 1;
	end	else if (num==16'd48973) begin
		AssumePrime = 1;
	end	else if (num==16'd48989) begin
		AssumePrime = 1;
	end	else if (num==16'd48991) begin
		AssumePrime = 1;
	end	else if (num==16'd49003) begin
		AssumePrime = 1;
	end	else if (num==16'd49009) begin
		AssumePrime = 1;
	end	else if (num==16'd49019) begin
		AssumePrime = 1;
	end	else if (num==16'd49031) begin
		AssumePrime = 1;
	end	else if (num==16'd49033) begin
		AssumePrime = 1;
	end	else if (num==16'd49037) begin
		AssumePrime = 1;
	end	else if (num==16'd49043) begin
		AssumePrime = 1;
	end	else if (num==16'd49057) begin
		AssumePrime = 1;
	end	else if (num==16'd49069) begin
		AssumePrime = 1;
	end	else if (num==16'd49081) begin
		AssumePrime = 1;
	end	else if (num==16'd49103) begin
		AssumePrime = 1;
	end	else if (num==16'd49109) begin
		AssumePrime = 1;
	end	else if (num==16'd49117) begin
		AssumePrime = 1;
	end	else if (num==16'd49121) begin
		AssumePrime = 1;
	end	else if (num==16'd49123) begin
		AssumePrime = 1;
	end	else if (num==16'd49139) begin
		AssumePrime = 1;
	end	else if (num==16'd49157) begin
		AssumePrime = 1;
	end	else if (num==16'd49169) begin
		AssumePrime = 1;
	end	else if (num==16'd49171) begin
		AssumePrime = 1;
	end	else if (num==16'd49177) begin
		AssumePrime = 1;
	end	else if (num==16'd49193) begin
		AssumePrime = 1;
	end	else if (num==16'd49199) begin
		AssumePrime = 1;
	end	else if (num==16'd49201) begin
		AssumePrime = 1;
	end	else if (num==16'd49207) begin
		AssumePrime = 1;
	end	else if (num==16'd49211) begin
		AssumePrime = 1;
	end	else if (num==16'd49223) begin
		AssumePrime = 1;
	end	else if (num==16'd49253) begin
		AssumePrime = 1;
	end	else if (num==16'd49261) begin
		AssumePrime = 1;
	end	else if (num==16'd49277) begin
		AssumePrime = 1;
	end	else if (num==16'd49279) begin
		AssumePrime = 1;
	end	else if (num==16'd49297) begin
		AssumePrime = 1;
	end	else if (num==16'd49307) begin
		AssumePrime = 1;
	end	else if (num==16'd49331) begin
		AssumePrime = 1;
	end	else if (num==16'd49333) begin
		AssumePrime = 1;
	end	else if (num==16'd49339) begin
		AssumePrime = 1;
	end	else if (num==16'd49363) begin
		AssumePrime = 1;
	end	else if (num==16'd49367) begin
		AssumePrime = 1;
	end	else if (num==16'd49369) begin
		AssumePrime = 1;
	end	else if (num==16'd49391) begin
		AssumePrime = 1;
	end	else if (num==16'd49393) begin
		AssumePrime = 1;
	end	else if (num==16'd49409) begin
		AssumePrime = 1;
	end	else if (num==16'd49411) begin
		AssumePrime = 1;
	end	else if (num==16'd49417) begin
		AssumePrime = 1;
	end	else if (num==16'd49429) begin
		AssumePrime = 1;
	end	else if (num==16'd49433) begin
		AssumePrime = 1;
	end	else if (num==16'd49451) begin
		AssumePrime = 1;
	end	else if (num==16'd49459) begin
		AssumePrime = 1;
	end	else if (num==16'd49463) begin
		AssumePrime = 1;
	end	else if (num==16'd49477) begin
		AssumePrime = 1;
	end	else if (num==16'd49481) begin
		AssumePrime = 1;
	end	else if (num==16'd49499) begin
		AssumePrime = 1;
	end	else if (num==16'd49523) begin
		AssumePrime = 1;
	end	else if (num==16'd49529) begin
		AssumePrime = 1;
	end	else if (num==16'd49531) begin
		AssumePrime = 1;
	end	else if (num==16'd49537) begin
		AssumePrime = 1;
	end	else if (num==16'd49547) begin
		AssumePrime = 1;
	end	else if (num==16'd49549) begin
		AssumePrime = 1;
	end	else if (num==16'd49559) begin
		AssumePrime = 1;
	end	else if (num==16'd49597) begin
		AssumePrime = 1;
	end	else if (num==16'd49603) begin
		AssumePrime = 1;
	end	else if (num==16'd49613) begin
		AssumePrime = 1;
	end	else if (num==16'd49627) begin
		AssumePrime = 1;
	end	else if (num==16'd49633) begin
		AssumePrime = 1;
	end	else if (num==16'd49639) begin
		AssumePrime = 1;
	end	else if (num==16'd49663) begin
		AssumePrime = 1;
	end	else if (num==16'd49667) begin
		AssumePrime = 1;
	end	else if (num==16'd49669) begin
		AssumePrime = 1;
	end	else if (num==16'd49681) begin
		AssumePrime = 1;
	end	else if (num==16'd49697) begin
		AssumePrime = 1;
	end	else if (num==16'd49711) begin
		AssumePrime = 1;
	end	else if (num==16'd49727) begin
		AssumePrime = 1;
	end	else if (num==16'd49739) begin
		AssumePrime = 1;
	end	else if (num==16'd49741) begin
		AssumePrime = 1;
	end	else if (num==16'd49747) begin
		AssumePrime = 1;
	end	else if (num==16'd49757) begin
		AssumePrime = 1;
	end	else if (num==16'd49783) begin
		AssumePrime = 1;
	end	else if (num==16'd49787) begin
		AssumePrime = 1;
	end	else if (num==16'd49789) begin
		AssumePrime = 1;
	end	else if (num==16'd49801) begin
		AssumePrime = 1;
	end	else if (num==16'd49807) begin
		AssumePrime = 1;
	end	else if (num==16'd49811) begin
		AssumePrime = 1;
	end	else if (num==16'd49823) begin
		AssumePrime = 1;
	end	else if (num==16'd49831) begin
		AssumePrime = 1;
	end	else if (num==16'd49843) begin
		AssumePrime = 1;
	end	else if (num==16'd49853) begin
		AssumePrime = 1;
	end	else if (num==16'd49871) begin
		AssumePrime = 1;
	end	else if (num==16'd49877) begin
		AssumePrime = 1;
	end	else if (num==16'd49891) begin
		AssumePrime = 1;
	end	else if (num==16'd49919) begin
		AssumePrime = 1;
	end	else if (num==16'd49921) begin
		AssumePrime = 1;
	end	else if (num==16'd49927) begin
		AssumePrime = 1;
	end	else if (num==16'd49937) begin
		AssumePrime = 1;
	end	else if (num==16'd49939) begin
		AssumePrime = 1;
	end	else if (num==16'd49943) begin
		AssumePrime = 1;
	end	else if (num==16'd49957) begin
		AssumePrime = 1;
	end	else if (num==16'd49991) begin
		AssumePrime = 1;
	end	else if (num==16'd49993) begin
		AssumePrime = 1;
	end	else if (num==16'd49999) begin
		AssumePrime = 1;
	end	else if (num==16'd50021) begin
		AssumePrime = 1;
	end	else if (num==16'd50023) begin
		AssumePrime = 1;
	end	else if (num==16'd50033) begin
		AssumePrime = 1;
	end	else if (num==16'd50047) begin
		AssumePrime = 1;
	end	else if (num==16'd50051) begin
		AssumePrime = 1;
	end	else if (num==16'd50053) begin
		AssumePrime = 1;
	end	else if (num==16'd50069) begin
		AssumePrime = 1;
	end	else if (num==16'd50077) begin
		AssumePrime = 1;
	end	else if (num==16'd50087) begin
		AssumePrime = 1;
	end	else if (num==16'd50093) begin
		AssumePrime = 1;
	end	else if (num==16'd50101) begin
		AssumePrime = 1;
	end	else if (num==16'd50111) begin
		AssumePrime = 1;
	end	else if (num==16'd50119) begin
		AssumePrime = 1;
	end	else if (num==16'd50123) begin
		AssumePrime = 1;
	end	else if (num==16'd50129) begin
		AssumePrime = 1;
	end	else if (num==16'd50131) begin
		AssumePrime = 1;
	end	else if (num==16'd50147) begin
		AssumePrime = 1;
	end	else if (num==16'd50153) begin
		AssumePrime = 1;
	end	else if (num==16'd50159) begin
		AssumePrime = 1;
	end	else if (num==16'd50177) begin
		AssumePrime = 1;
	end	else if (num==16'd50207) begin
		AssumePrime = 1;
	end	else if (num==16'd50221) begin
		AssumePrime = 1;
	end	else if (num==16'd50227) begin
		AssumePrime = 1;
	end	else if (num==16'd50231) begin
		AssumePrime = 1;
	end	else if (num==16'd50261) begin
		AssumePrime = 1;
	end	else if (num==16'd50263) begin
		AssumePrime = 1;
	end	else if (num==16'd50273) begin
		AssumePrime = 1;
	end	else if (num==16'd50287) begin
		AssumePrime = 1;
	end	else if (num==16'd50291) begin
		AssumePrime = 1;
	end	else if (num==16'd50311) begin
		AssumePrime = 1;
	end	else if (num==16'd50321) begin
		AssumePrime = 1;
	end	else if (num==16'd50329) begin
		AssumePrime = 1;
	end	else if (num==16'd50333) begin
		AssumePrime = 1;
	end	else if (num==16'd50341) begin
		AssumePrime = 1;
	end	else if (num==16'd50359) begin
		AssumePrime = 1;
	end	else if (num==16'd50363) begin
		AssumePrime = 1;
	end	else if (num==16'd50377) begin
		AssumePrime = 1;
	end	else if (num==16'd50383) begin
		AssumePrime = 1;
	end	else if (num==16'd50387) begin
		AssumePrime = 1;
	end	else if (num==16'd50411) begin
		AssumePrime = 1;
	end	else if (num==16'd50417) begin
		AssumePrime = 1;
	end	else if (num==16'd50423) begin
		AssumePrime = 1;
	end	else if (num==16'd50441) begin
		AssumePrime = 1;
	end	else if (num==16'd50459) begin
		AssumePrime = 1;
	end	else if (num==16'd50461) begin
		AssumePrime = 1;
	end	else if (num==16'd50497) begin
		AssumePrime = 1;
	end	else if (num==16'd50503) begin
		AssumePrime = 1;
	end	else if (num==16'd50513) begin
		AssumePrime = 1;
	end	else if (num==16'd50527) begin
		AssumePrime = 1;
	end	else if (num==16'd50539) begin
		AssumePrime = 1;
	end	else if (num==16'd50543) begin
		AssumePrime = 1;
	end	else if (num==16'd50549) begin
		AssumePrime = 1;
	end	else if (num==16'd50551) begin
		AssumePrime = 1;
	end	else if (num==16'd50581) begin
		AssumePrime = 1;
	end	else if (num==16'd50587) begin
		AssumePrime = 1;
	end	else if (num==16'd50591) begin
		AssumePrime = 1;
	end	else if (num==16'd50593) begin
		AssumePrime = 1;
	end	else if (num==16'd50599) begin
		AssumePrime = 1;
	end	else if (num==16'd50627) begin
		AssumePrime = 1;
	end	else if (num==16'd50647) begin
		AssumePrime = 1;
	end	else if (num==16'd50651) begin
		AssumePrime = 1;
	end	else if (num==16'd50671) begin
		AssumePrime = 1;
	end	else if (num==16'd50683) begin
		AssumePrime = 1;
	end	else if (num==16'd50707) begin
		AssumePrime = 1;
	end	else if (num==16'd50723) begin
		AssumePrime = 1;
	end	else if (num==16'd50741) begin
		AssumePrime = 1;
	end	else if (num==16'd50753) begin
		AssumePrime = 1;
	end	else if (num==16'd50767) begin
		AssumePrime = 1;
	end	else if (num==16'd50773) begin
		AssumePrime = 1;
	end	else if (num==16'd50777) begin
		AssumePrime = 1;
	end	else if (num==16'd50789) begin
		AssumePrime = 1;
	end	else if (num==16'd50821) begin
		AssumePrime = 1;
	end	else if (num==16'd50833) begin
		AssumePrime = 1;
	end	else if (num==16'd50839) begin
		AssumePrime = 1;
	end	else if (num==16'd50849) begin
		AssumePrime = 1;
	end	else if (num==16'd50857) begin
		AssumePrime = 1;
	end	else if (num==16'd50867) begin
		AssumePrime = 1;
	end	else if (num==16'd50873) begin
		AssumePrime = 1;
	end	else if (num==16'd50891) begin
		AssumePrime = 1;
	end	else if (num==16'd50893) begin
		AssumePrime = 1;
	end	else if (num==16'd50909) begin
		AssumePrime = 1;
	end	else if (num==16'd50923) begin
		AssumePrime = 1;
	end	else if (num==16'd50929) begin
		AssumePrime = 1;
	end	else if (num==16'd50951) begin
		AssumePrime = 1;
	end	else if (num==16'd50957) begin
		AssumePrime = 1;
	end	else if (num==16'd50969) begin
		AssumePrime = 1;
	end	else if (num==16'd50971) begin
		AssumePrime = 1;
	end	else if (num==16'd50989) begin
		AssumePrime = 1;
	end	else if (num==16'd50993) begin
		AssumePrime = 1;
	end	else if (num==16'd51001) begin
		AssumePrime = 1;
	end	else if (num==16'd51031) begin
		AssumePrime = 1;
	end	else if (num==16'd51043) begin
		AssumePrime = 1;
	end	else if (num==16'd51047) begin
		AssumePrime = 1;
	end	else if (num==16'd51059) begin
		AssumePrime = 1;
	end	else if (num==16'd51061) begin
		AssumePrime = 1;
	end	else if (num==16'd51071) begin
		AssumePrime = 1;
	end	else if (num==16'd51109) begin
		AssumePrime = 1;
	end	else if (num==16'd51131) begin
		AssumePrime = 1;
	end	else if (num==16'd51133) begin
		AssumePrime = 1;
	end	else if (num==16'd51137) begin
		AssumePrime = 1;
	end	else if (num==16'd51151) begin
		AssumePrime = 1;
	end	else if (num==16'd51157) begin
		AssumePrime = 1;
	end	else if (num==16'd51169) begin
		AssumePrime = 1;
	end	else if (num==16'd51193) begin
		AssumePrime = 1;
	end	else if (num==16'd51197) begin
		AssumePrime = 1;
	end	else if (num==16'd51199) begin
		AssumePrime = 1;
	end	else if (num==16'd51203) begin
		AssumePrime = 1;
	end	else if (num==16'd51217) begin
		AssumePrime = 1;
	end	else if (num==16'd51229) begin
		AssumePrime = 1;
	end	else if (num==16'd51239) begin
		AssumePrime = 1;
	end	else if (num==16'd51241) begin
		AssumePrime = 1;
	end	else if (num==16'd51257) begin
		AssumePrime = 1;
	end	else if (num==16'd51263) begin
		AssumePrime = 1;
	end	else if (num==16'd51283) begin
		AssumePrime = 1;
	end	else if (num==16'd51287) begin
		AssumePrime = 1;
	end	else if (num==16'd51307) begin
		AssumePrime = 1;
	end	else if (num==16'd51329) begin
		AssumePrime = 1;
	end	else if (num==16'd51341) begin
		AssumePrime = 1;
	end	else if (num==16'd51343) begin
		AssumePrime = 1;
	end	else if (num==16'd51347) begin
		AssumePrime = 1;
	end	else if (num==16'd51349) begin
		AssumePrime = 1;
	end	else if (num==16'd51361) begin
		AssumePrime = 1;
	end	else if (num==16'd51383) begin
		AssumePrime = 1;
	end	else if (num==16'd51407) begin
		AssumePrime = 1;
	end	else if (num==16'd51413) begin
		AssumePrime = 1;
	end	else if (num==16'd51419) begin
		AssumePrime = 1;
	end	else if (num==16'd51421) begin
		AssumePrime = 1;
	end	else if (num==16'd51427) begin
		AssumePrime = 1;
	end	else if (num==16'd51431) begin
		AssumePrime = 1;
	end	else if (num==16'd51437) begin
		AssumePrime = 1;
	end	else if (num==16'd51439) begin
		AssumePrime = 1;
	end	else if (num==16'd51449) begin
		AssumePrime = 1;
	end	else if (num==16'd51461) begin
		AssumePrime = 1;
	end	else if (num==16'd51473) begin
		AssumePrime = 1;
	end	else if (num==16'd51479) begin
		AssumePrime = 1;
	end	else if (num==16'd51481) begin
		AssumePrime = 1;
	end	else if (num==16'd51487) begin
		AssumePrime = 1;
	end	else if (num==16'd51503) begin
		AssumePrime = 1;
	end	else if (num==16'd51511) begin
		AssumePrime = 1;
	end	else if (num==16'd51517) begin
		AssumePrime = 1;
	end	else if (num==16'd51521) begin
		AssumePrime = 1;
	end	else if (num==16'd51539) begin
		AssumePrime = 1;
	end	else if (num==16'd51551) begin
		AssumePrime = 1;
	end	else if (num==16'd51563) begin
		AssumePrime = 1;
	end	else if (num==16'd51577) begin
		AssumePrime = 1;
	end	else if (num==16'd51581) begin
		AssumePrime = 1;
	end	else if (num==16'd51593) begin
		AssumePrime = 1;
	end	else if (num==16'd51599) begin
		AssumePrime = 1;
	end	else if (num==16'd51607) begin
		AssumePrime = 1;
	end	else if (num==16'd51613) begin
		AssumePrime = 1;
	end	else if (num==16'd51631) begin
		AssumePrime = 1;
	end	else if (num==16'd51637) begin
		AssumePrime = 1;
	end	else if (num==16'd51647) begin
		AssumePrime = 1;
	end	else if (num==16'd51659) begin
		AssumePrime = 1;
	end	else if (num==16'd51673) begin
		AssumePrime = 1;
	end	else if (num==16'd51679) begin
		AssumePrime = 1;
	end	else if (num==16'd51683) begin
		AssumePrime = 1;
	end	else if (num==16'd51691) begin
		AssumePrime = 1;
	end	else if (num==16'd51713) begin
		AssumePrime = 1;
	end	else if (num==16'd51719) begin
		AssumePrime = 1;
	end	else if (num==16'd51721) begin
		AssumePrime = 1;
	end	else if (num==16'd51749) begin
		AssumePrime = 1;
	end	else if (num==16'd51767) begin
		AssumePrime = 1;
	end	else if (num==16'd51769) begin
		AssumePrime = 1;
	end	else if (num==16'd51787) begin
		AssumePrime = 1;
	end	else if (num==16'd51797) begin
		AssumePrime = 1;
	end	else if (num==16'd51803) begin
		AssumePrime = 1;
	end	else if (num==16'd51817) begin
		AssumePrime = 1;
	end	else if (num==16'd51827) begin
		AssumePrime = 1;
	end	else if (num==16'd51829) begin
		AssumePrime = 1;
	end	else if (num==16'd51839) begin
		AssumePrime = 1;
	end	else if (num==16'd51853) begin
		AssumePrime = 1;
	end	else if (num==16'd51859) begin
		AssumePrime = 1;
	end	else if (num==16'd51869) begin
		AssumePrime = 1;
	end	else if (num==16'd51871) begin
		AssumePrime = 1;
	end	else if (num==16'd51893) begin
		AssumePrime = 1;
	end	else if (num==16'd51899) begin
		AssumePrime = 1;
	end	else if (num==16'd51907) begin
		AssumePrime = 1;
	end	else if (num==16'd51913) begin
		AssumePrime = 1;
	end	else if (num==16'd51929) begin
		AssumePrime = 1;
	end	else if (num==16'd51941) begin
		AssumePrime = 1;
	end	else if (num==16'd51949) begin
		AssumePrime = 1;
	end	else if (num==16'd51971) begin
		AssumePrime = 1;
	end	else if (num==16'd51973) begin
		AssumePrime = 1;
	end	else if (num==16'd51977) begin
		AssumePrime = 1;
	end	else if (num==16'd51991) begin
		AssumePrime = 1;
	end	else if (num==16'd52009) begin
		AssumePrime = 1;
	end	else if (num==16'd52021) begin
		AssumePrime = 1;
	end	else if (num==16'd52027) begin
		AssumePrime = 1;
	end	else if (num==16'd52051) begin
		AssumePrime = 1;
	end	else if (num==16'd52057) begin
		AssumePrime = 1;
	end	else if (num==16'd52067) begin
		AssumePrime = 1;
	end	else if (num==16'd52069) begin
		AssumePrime = 1;
	end	else if (num==16'd52081) begin
		AssumePrime = 1;
	end	else if (num==16'd52103) begin
		AssumePrime = 1;
	end	else if (num==16'd52121) begin
		AssumePrime = 1;
	end	else if (num==16'd52127) begin
		AssumePrime = 1;
	end	else if (num==16'd52147) begin
		AssumePrime = 1;
	end	else if (num==16'd52153) begin
		AssumePrime = 1;
	end	else if (num==16'd52163) begin
		AssumePrime = 1;
	end	else if (num==16'd52177) begin
		AssumePrime = 1;
	end	else if (num==16'd52181) begin
		AssumePrime = 1;
	end	else if (num==16'd52183) begin
		AssumePrime = 1;
	end	else if (num==16'd52189) begin
		AssumePrime = 1;
	end	else if (num==16'd52201) begin
		AssumePrime = 1;
	end	else if (num==16'd52223) begin
		AssumePrime = 1;
	end	else if (num==16'd52237) begin
		AssumePrime = 1;
	end	else if (num==16'd52249) begin
		AssumePrime = 1;
	end	else if (num==16'd52253) begin
		AssumePrime = 1;
	end	else if (num==16'd52259) begin
		AssumePrime = 1;
	end	else if (num==16'd52267) begin
		AssumePrime = 1;
	end	else if (num==16'd52289) begin
		AssumePrime = 1;
	end	else if (num==16'd52291) begin
		AssumePrime = 1;
	end	else if (num==16'd52301) begin
		AssumePrime = 1;
	end	else if (num==16'd52313) begin
		AssumePrime = 1;
	end	else if (num==16'd52321) begin
		AssumePrime = 1;
	end	else if (num==16'd52361) begin
		AssumePrime = 1;
	end	else if (num==16'd52363) begin
		AssumePrime = 1;
	end	else if (num==16'd52369) begin
		AssumePrime = 1;
	end	else if (num==16'd52379) begin
		AssumePrime = 1;
	end	else if (num==16'd52387) begin
		AssumePrime = 1;
	end	else if (num==16'd52391) begin
		AssumePrime = 1;
	end	else if (num==16'd52433) begin
		AssumePrime = 1;
	end	else if (num==16'd52453) begin
		AssumePrime = 1;
	end	else if (num==16'd52457) begin
		AssumePrime = 1;
	end	else if (num==16'd52489) begin
		AssumePrime = 1;
	end	else if (num==16'd52501) begin
		AssumePrime = 1;
	end	else if (num==16'd52511) begin
		AssumePrime = 1;
	end	else if (num==16'd52517) begin
		AssumePrime = 1;
	end	else if (num==16'd52529) begin
		AssumePrime = 1;
	end	else if (num==16'd52541) begin
		AssumePrime = 1;
	end	else if (num==16'd52543) begin
		AssumePrime = 1;
	end	else if (num==16'd52553) begin
		AssumePrime = 1;
	end	else if (num==16'd52561) begin
		AssumePrime = 1;
	end	else if (num==16'd52567) begin
		AssumePrime = 1;
	end	else if (num==16'd52571) begin
		AssumePrime = 1;
	end	else if (num==16'd52579) begin
		AssumePrime = 1;
	end	else if (num==16'd52583) begin
		AssumePrime = 1;
	end	else if (num==16'd52609) begin
		AssumePrime = 1;
	end	else if (num==16'd52627) begin
		AssumePrime = 1;
	end	else if (num==16'd52631) begin
		AssumePrime = 1;
	end	else if (num==16'd52639) begin
		AssumePrime = 1;
	end	else if (num==16'd52667) begin
		AssumePrime = 1;
	end	else if (num==16'd52673) begin
		AssumePrime = 1;
	end	else if (num==16'd52691) begin
		AssumePrime = 1;
	end	else if (num==16'd52697) begin
		AssumePrime = 1;
	end	else if (num==16'd52709) begin
		AssumePrime = 1;
	end	else if (num==16'd52711) begin
		AssumePrime = 1;
	end	else if (num==16'd52721) begin
		AssumePrime = 1;
	end	else if (num==16'd52727) begin
		AssumePrime = 1;
	end	else if (num==16'd52733) begin
		AssumePrime = 1;
	end	else if (num==16'd52747) begin
		AssumePrime = 1;
	end	else if (num==16'd52757) begin
		AssumePrime = 1;
	end	else if (num==16'd52769) begin
		AssumePrime = 1;
	end	else if (num==16'd52783) begin
		AssumePrime = 1;
	end	else if (num==16'd52807) begin
		AssumePrime = 1;
	end	else if (num==16'd52813) begin
		AssumePrime = 1;
	end	else if (num==16'd52817) begin
		AssumePrime = 1;
	end	else if (num==16'd52837) begin
		AssumePrime = 1;
	end	else if (num==16'd52859) begin
		AssumePrime = 1;
	end	else if (num==16'd52861) begin
		AssumePrime = 1;
	end	else if (num==16'd52879) begin
		AssumePrime = 1;
	end	else if (num==16'd52883) begin
		AssumePrime = 1;
	end	else if (num==16'd52889) begin
		AssumePrime = 1;
	end	else if (num==16'd52901) begin
		AssumePrime = 1;
	end	else if (num==16'd52903) begin
		AssumePrime = 1;
	end	else if (num==16'd52919) begin
		AssumePrime = 1;
	end	else if (num==16'd52937) begin
		AssumePrime = 1;
	end	else if (num==16'd52951) begin
		AssumePrime = 1;
	end	else if (num==16'd52957) begin
		AssumePrime = 1;
	end	else if (num==16'd52963) begin
		AssumePrime = 1;
	end	else if (num==16'd52967) begin
		AssumePrime = 1;
	end	else if (num==16'd52973) begin
		AssumePrime = 1;
	end	else if (num==16'd52981) begin
		AssumePrime = 1;
	end	else if (num==16'd52999) begin
		AssumePrime = 1;
	end	else if (num==16'd53003) begin
		AssumePrime = 1;
	end	else if (num==16'd53017) begin
		AssumePrime = 1;
	end	else if (num==16'd53047) begin
		AssumePrime = 1;
	end	else if (num==16'd53051) begin
		AssumePrime = 1;
	end	else if (num==16'd53069) begin
		AssumePrime = 1;
	end	else if (num==16'd53077) begin
		AssumePrime = 1;
	end	else if (num==16'd53087) begin
		AssumePrime = 1;
	end	else if (num==16'd53089) begin
		AssumePrime = 1;
	end	else if (num==16'd53093) begin
		AssumePrime = 1;
	end	else if (num==16'd53101) begin
		AssumePrime = 1;
	end	else if (num==16'd53113) begin
		AssumePrime = 1;
	end	else if (num==16'd53117) begin
		AssumePrime = 1;
	end	else if (num==16'd53129) begin
		AssumePrime = 1;
	end	else if (num==16'd53147) begin
		AssumePrime = 1;
	end	else if (num==16'd53149) begin
		AssumePrime = 1;
	end	else if (num==16'd53161) begin
		AssumePrime = 1;
	end	else if (num==16'd53171) begin
		AssumePrime = 1;
	end	else if (num==16'd53173) begin
		AssumePrime = 1;
	end	else if (num==16'd53189) begin
		AssumePrime = 1;
	end	else if (num==16'd53197) begin
		AssumePrime = 1;
	end	else if (num==16'd53201) begin
		AssumePrime = 1;
	end	else if (num==16'd53231) begin
		AssumePrime = 1;
	end	else if (num==16'd53233) begin
		AssumePrime = 1;
	end	else if (num==16'd53239) begin
		AssumePrime = 1;
	end	else if (num==16'd53267) begin
		AssumePrime = 1;
	end	else if (num==16'd53269) begin
		AssumePrime = 1;
	end	else if (num==16'd53279) begin
		AssumePrime = 1;
	end	else if (num==16'd53281) begin
		AssumePrime = 1;
	end	else if (num==16'd53299) begin
		AssumePrime = 1;
	end	else if (num==16'd53309) begin
		AssumePrime = 1;
	end	else if (num==16'd53323) begin
		AssumePrime = 1;
	end	else if (num==16'd53327) begin
		AssumePrime = 1;
	end	else if (num==16'd53353) begin
		AssumePrime = 1;
	end	else if (num==16'd53359) begin
		AssumePrime = 1;
	end	else if (num==16'd53377) begin
		AssumePrime = 1;
	end	else if (num==16'd53381) begin
		AssumePrime = 1;
	end	else if (num==16'd53401) begin
		AssumePrime = 1;
	end	else if (num==16'd53407) begin
		AssumePrime = 1;
	end	else if (num==16'd53411) begin
		AssumePrime = 1;
	end	else if (num==16'd53419) begin
		AssumePrime = 1;
	end	else if (num==16'd53437) begin
		AssumePrime = 1;
	end	else if (num==16'd53441) begin
		AssumePrime = 1;
	end	else if (num==16'd53453) begin
		AssumePrime = 1;
	end	else if (num==16'd53479) begin
		AssumePrime = 1;
	end	else if (num==16'd53503) begin
		AssumePrime = 1;
	end	else if (num==16'd53507) begin
		AssumePrime = 1;
	end	else if (num==16'd53527) begin
		AssumePrime = 1;
	end	else if (num==16'd53549) begin
		AssumePrime = 1;
	end	else if (num==16'd53551) begin
		AssumePrime = 1;
	end	else if (num==16'd53569) begin
		AssumePrime = 1;
	end	else if (num==16'd53591) begin
		AssumePrime = 1;
	end	else if (num==16'd53593) begin
		AssumePrime = 1;
	end	else if (num==16'd53597) begin
		AssumePrime = 1;
	end	else if (num==16'd53609) begin
		AssumePrime = 1;
	end	else if (num==16'd53611) begin
		AssumePrime = 1;
	end	else if (num==16'd53617) begin
		AssumePrime = 1;
	end	else if (num==16'd53623) begin
		AssumePrime = 1;
	end	else if (num==16'd53629) begin
		AssumePrime = 1;
	end	else if (num==16'd53633) begin
		AssumePrime = 1;
	end	else if (num==16'd53639) begin
		AssumePrime = 1;
	end	else if (num==16'd53653) begin
		AssumePrime = 1;
	end	else if (num==16'd53657) begin
		AssumePrime = 1;
	end	else if (num==16'd53681) begin
		AssumePrime = 1;
	end	else if (num==16'd53693) begin
		AssumePrime = 1;
	end	else if (num==16'd53699) begin
		AssumePrime = 1;
	end	else if (num==16'd53717) begin
		AssumePrime = 1;
	end	else if (num==16'd53719) begin
		AssumePrime = 1;
	end	else if (num==16'd53731) begin
		AssumePrime = 1;
	end	else if (num==16'd53759) begin
		AssumePrime = 1;
	end	else if (num==16'd53773) begin
		AssumePrime = 1;
	end	else if (num==16'd53777) begin
		AssumePrime = 1;
	end	else if (num==16'd53783) begin
		AssumePrime = 1;
	end	else if (num==16'd53791) begin
		AssumePrime = 1;
	end	else if (num==16'd53813) begin
		AssumePrime = 1;
	end	else if (num==16'd53819) begin
		AssumePrime = 1;
	end	else if (num==16'd53831) begin
		AssumePrime = 1;
	end	else if (num==16'd53849) begin
		AssumePrime = 1;
	end	else if (num==16'd53857) begin
		AssumePrime = 1;
	end	else if (num==16'd53861) begin
		AssumePrime = 1;
	end	else if (num==16'd53881) begin
		AssumePrime = 1;
	end	else if (num==16'd53887) begin
		AssumePrime = 1;
	end	else if (num==16'd53891) begin
		AssumePrime = 1;
	end	else if (num==16'd53897) begin
		AssumePrime = 1;
	end	else if (num==16'd53899) begin
		AssumePrime = 1;
	end	else if (num==16'd53917) begin
		AssumePrime = 1;
	end	else if (num==16'd53923) begin
		AssumePrime = 1;
	end	else if (num==16'd53927) begin
		AssumePrime = 1;
	end	else if (num==16'd53939) begin
		AssumePrime = 1;
	end	else if (num==16'd53951) begin
		AssumePrime = 1;
	end	else if (num==16'd53959) begin
		AssumePrime = 1;
	end	else if (num==16'd53987) begin
		AssumePrime = 1;
	end	else if (num==16'd53993) begin
		AssumePrime = 1;
	end	else if (num==16'd54001) begin
		AssumePrime = 1;
	end	else if (num==16'd54011) begin
		AssumePrime = 1;
	end	else if (num==16'd54013) begin
		AssumePrime = 1;
	end	else if (num==16'd54037) begin
		AssumePrime = 1;
	end	else if (num==16'd54049) begin
		AssumePrime = 1;
	end	else if (num==16'd54059) begin
		AssumePrime = 1;
	end	else if (num==16'd54083) begin
		AssumePrime = 1;
	end	else if (num==16'd54091) begin
		AssumePrime = 1;
	end	else if (num==16'd54101) begin
		AssumePrime = 1;
	end	else if (num==16'd54121) begin
		AssumePrime = 1;
	end	else if (num==16'd54133) begin
		AssumePrime = 1;
	end	else if (num==16'd54139) begin
		AssumePrime = 1;
	end	else if (num==16'd54151) begin
		AssumePrime = 1;
	end	else if (num==16'd54163) begin
		AssumePrime = 1;
	end	else if (num==16'd54167) begin
		AssumePrime = 1;
	end	else if (num==16'd54181) begin
		AssumePrime = 1;
	end	else if (num==16'd54193) begin
		AssumePrime = 1;
	end	else if (num==16'd54217) begin
		AssumePrime = 1;
	end	else if (num==16'd54251) begin
		AssumePrime = 1;
	end	else if (num==16'd54269) begin
		AssumePrime = 1;
	end	else if (num==16'd54277) begin
		AssumePrime = 1;
	end	else if (num==16'd54287) begin
		AssumePrime = 1;
	end	else if (num==16'd54293) begin
		AssumePrime = 1;
	end	else if (num==16'd54311) begin
		AssumePrime = 1;
	end	else if (num==16'd54319) begin
		AssumePrime = 1;
	end	else if (num==16'd54323) begin
		AssumePrime = 1;
	end	else if (num==16'd54331) begin
		AssumePrime = 1;
	end	else if (num==16'd54347) begin
		AssumePrime = 1;
	end	else if (num==16'd54361) begin
		AssumePrime = 1;
	end	else if (num==16'd54367) begin
		AssumePrime = 1;
	end	else if (num==16'd54371) begin
		AssumePrime = 1;
	end	else if (num==16'd54377) begin
		AssumePrime = 1;
	end	else if (num==16'd54401) begin
		AssumePrime = 1;
	end	else if (num==16'd54403) begin
		AssumePrime = 1;
	end	else if (num==16'd54409) begin
		AssumePrime = 1;
	end	else if (num==16'd54413) begin
		AssumePrime = 1;
	end	else if (num==16'd54419) begin
		AssumePrime = 1;
	end	else if (num==16'd54421) begin
		AssumePrime = 1;
	end	else if (num==16'd54437) begin
		AssumePrime = 1;
	end	else if (num==16'd54443) begin
		AssumePrime = 1;
	end	else if (num==16'd54449) begin
		AssumePrime = 1;
	end	else if (num==16'd54469) begin
		AssumePrime = 1;
	end	else if (num==16'd54493) begin
		AssumePrime = 1;
	end	else if (num==16'd54497) begin
		AssumePrime = 1;
	end	else if (num==16'd54499) begin
		AssumePrime = 1;
	end	else if (num==16'd54503) begin
		AssumePrime = 1;
	end	else if (num==16'd54517) begin
		AssumePrime = 1;
	end	else if (num==16'd54521) begin
		AssumePrime = 1;
	end	else if (num==16'd54539) begin
		AssumePrime = 1;
	end	else if (num==16'd54541) begin
		AssumePrime = 1;
	end	else if (num==16'd54547) begin
		AssumePrime = 1;
	end	else if (num==16'd54559) begin
		AssumePrime = 1;
	end	else if (num==16'd54563) begin
		AssumePrime = 1;
	end	else if (num==16'd54577) begin
		AssumePrime = 1;
	end	else if (num==16'd54581) begin
		AssumePrime = 1;
	end	else if (num==16'd54583) begin
		AssumePrime = 1;
	end	else if (num==16'd54601) begin
		AssumePrime = 1;
	end	else if (num==16'd54617) begin
		AssumePrime = 1;
	end	else if (num==16'd54623) begin
		AssumePrime = 1;
	end	else if (num==16'd54629) begin
		AssumePrime = 1;
	end	else if (num==16'd54631) begin
		AssumePrime = 1;
	end	else if (num==16'd54647) begin
		AssumePrime = 1;
	end	else if (num==16'd54667) begin
		AssumePrime = 1;
	end	else if (num==16'd54673) begin
		AssumePrime = 1;
	end	else if (num==16'd54679) begin
		AssumePrime = 1;
	end	else if (num==16'd54709) begin
		AssumePrime = 1;
	end	else if (num==16'd54713) begin
		AssumePrime = 1;
	end	else if (num==16'd54721) begin
		AssumePrime = 1;
	end	else if (num==16'd54727) begin
		AssumePrime = 1;
	end	else if (num==16'd54751) begin
		AssumePrime = 1;
	end	else if (num==16'd54767) begin
		AssumePrime = 1;
	end	else if (num==16'd54773) begin
		AssumePrime = 1;
	end	else if (num==16'd54779) begin
		AssumePrime = 1;
	end	else if (num==16'd54787) begin
		AssumePrime = 1;
	end	else if (num==16'd54799) begin
		AssumePrime = 1;
	end	else if (num==16'd54829) begin
		AssumePrime = 1;
	end	else if (num==16'd54833) begin
		AssumePrime = 1;
	end	else if (num==16'd54851) begin
		AssumePrime = 1;
	end	else if (num==16'd54869) begin
		AssumePrime = 1;
	end	else if (num==16'd54877) begin
		AssumePrime = 1;
	end	else if (num==16'd54881) begin
		AssumePrime = 1;
	end	else if (num==16'd54907) begin
		AssumePrime = 1;
	end	else if (num==16'd54917) begin
		AssumePrime = 1;
	end	else if (num==16'd54919) begin
		AssumePrime = 1;
	end	else if (num==16'd54941) begin
		AssumePrime = 1;
	end	else if (num==16'd54949) begin
		AssumePrime = 1;
	end	else if (num==16'd54959) begin
		AssumePrime = 1;
	end	else if (num==16'd54973) begin
		AssumePrime = 1;
	end	else if (num==16'd54979) begin
		AssumePrime = 1;
	end	else if (num==16'd54983) begin
		AssumePrime = 1;
	end	else if (num==16'd55001) begin
		AssumePrime = 1;
	end	else if (num==16'd55009) begin
		AssumePrime = 1;
	end	else if (num==16'd55021) begin
		AssumePrime = 1;
	end	else if (num==16'd55049) begin
		AssumePrime = 1;
	end	else if (num==16'd55051) begin
		AssumePrime = 1;
	end	else if (num==16'd55057) begin
		AssumePrime = 1;
	end	else if (num==16'd55061) begin
		AssumePrime = 1;
	end	else if (num==16'd55073) begin
		AssumePrime = 1;
	end	else if (num==16'd55079) begin
		AssumePrime = 1;
	end	else if (num==16'd55103) begin
		AssumePrime = 1;
	end	else if (num==16'd55109) begin
		AssumePrime = 1;
	end	else if (num==16'd55117) begin
		AssumePrime = 1;
	end	else if (num==16'd55127) begin
		AssumePrime = 1;
	end	else if (num==16'd55147) begin
		AssumePrime = 1;
	end	else if (num==16'd55163) begin
		AssumePrime = 1;
	end	else if (num==16'd55171) begin
		AssumePrime = 1;
	end	else if (num==16'd55201) begin
		AssumePrime = 1;
	end	else if (num==16'd55207) begin
		AssumePrime = 1;
	end	else if (num==16'd55213) begin
		AssumePrime = 1;
	end	else if (num==16'd55217) begin
		AssumePrime = 1;
	end	else if (num==16'd55219) begin
		AssumePrime = 1;
	end	else if (num==16'd55229) begin
		AssumePrime = 1;
	end	else if (num==16'd55243) begin
		AssumePrime = 1;
	end	else if (num==16'd55249) begin
		AssumePrime = 1;
	end	else if (num==16'd55259) begin
		AssumePrime = 1;
	end	else if (num==16'd55291) begin
		AssumePrime = 1;
	end	else if (num==16'd55313) begin
		AssumePrime = 1;
	end	else if (num==16'd55331) begin
		AssumePrime = 1;
	end	else if (num==16'd55333) begin
		AssumePrime = 1;
	end	else if (num==16'd55337) begin
		AssumePrime = 1;
	end	else if (num==16'd55339) begin
		AssumePrime = 1;
	end	else if (num==16'd55343) begin
		AssumePrime = 1;
	end	else if (num==16'd55351) begin
		AssumePrime = 1;
	end	else if (num==16'd55373) begin
		AssumePrime = 1;
	end	else if (num==16'd55381) begin
		AssumePrime = 1;
	end	else if (num==16'd55399) begin
		AssumePrime = 1;
	end	else if (num==16'd55411) begin
		AssumePrime = 1;
	end	else if (num==16'd55439) begin
		AssumePrime = 1;
	end	else if (num==16'd55441) begin
		AssumePrime = 1;
	end	else if (num==16'd55457) begin
		AssumePrime = 1;
	end	else if (num==16'd55469) begin
		AssumePrime = 1;
	end	else if (num==16'd55487) begin
		AssumePrime = 1;
	end	else if (num==16'd55501) begin
		AssumePrime = 1;
	end	else if (num==16'd55511) begin
		AssumePrime = 1;
	end	else if (num==16'd55529) begin
		AssumePrime = 1;
	end	else if (num==16'd55541) begin
		AssumePrime = 1;
	end	else if (num==16'd55547) begin
		AssumePrime = 1;
	end	else if (num==16'd55579) begin
		AssumePrime = 1;
	end	else if (num==16'd55589) begin
		AssumePrime = 1;
	end	else if (num==16'd55603) begin
		AssumePrime = 1;
	end	else if (num==16'd55609) begin
		AssumePrime = 1;
	end	else if (num==16'd55619) begin
		AssumePrime = 1;
	end	else if (num==16'd55621) begin
		AssumePrime = 1;
	end	else if (num==16'd55631) begin
		AssumePrime = 1;
	end	else if (num==16'd55633) begin
		AssumePrime = 1;
	end	else if (num==16'd55639) begin
		AssumePrime = 1;
	end	else if (num==16'd55661) begin
		AssumePrime = 1;
	end	else if (num==16'd55663) begin
		AssumePrime = 1;
	end	else if (num==16'd55667) begin
		AssumePrime = 1;
	end	else if (num==16'd55673) begin
		AssumePrime = 1;
	end	else if (num==16'd55681) begin
		AssumePrime = 1;
	end	else if (num==16'd55691) begin
		AssumePrime = 1;
	end	else if (num==16'd55697) begin
		AssumePrime = 1;
	end	else if (num==16'd55711) begin
		AssumePrime = 1;
	end	else if (num==16'd55717) begin
		AssumePrime = 1;
	end	else if (num==16'd55721) begin
		AssumePrime = 1;
	end	else if (num==16'd55733) begin
		AssumePrime = 1;
	end	else if (num==16'd55763) begin
		AssumePrime = 1;
	end	else if (num==16'd55787) begin
		AssumePrime = 1;
	end	else if (num==16'd55793) begin
		AssumePrime = 1;
	end	else if (num==16'd55799) begin
		AssumePrime = 1;
	end	else if (num==16'd55807) begin
		AssumePrime = 1;
	end	else if (num==16'd55813) begin
		AssumePrime = 1;
	end	else if (num==16'd55817) begin
		AssumePrime = 1;
	end	else if (num==16'd55819) begin
		AssumePrime = 1;
	end	else if (num==16'd55823) begin
		AssumePrime = 1;
	end	else if (num==16'd55829) begin
		AssumePrime = 1;
	end	else if (num==16'd55837) begin
		AssumePrime = 1;
	end	else if (num==16'd55843) begin
		AssumePrime = 1;
	end	else if (num==16'd55849) begin
		AssumePrime = 1;
	end	else if (num==16'd55871) begin
		AssumePrime = 1;
	end	else if (num==16'd55889) begin
		AssumePrime = 1;
	end	else if (num==16'd55897) begin
		AssumePrime = 1;
	end	else if (num==16'd55901) begin
		AssumePrime = 1;
	end	else if (num==16'd55903) begin
		AssumePrime = 1;
	end	else if (num==16'd55921) begin
		AssumePrime = 1;
	end	else if (num==16'd55927) begin
		AssumePrime = 1;
	end	else if (num==16'd55931) begin
		AssumePrime = 1;
	end	else if (num==16'd55933) begin
		AssumePrime = 1;
	end	else if (num==16'd55949) begin
		AssumePrime = 1;
	end	else if (num==16'd55967) begin
		AssumePrime = 1;
	end	else if (num==16'd55987) begin
		AssumePrime = 1;
	end	else if (num==16'd55997) begin
		AssumePrime = 1;
	end	else if (num==16'd56003) begin
		AssumePrime = 1;
	end	else if (num==16'd56009) begin
		AssumePrime = 1;
	end	else if (num==16'd56039) begin
		AssumePrime = 1;
	end	else if (num==16'd56041) begin
		AssumePrime = 1;
	end	else if (num==16'd56053) begin
		AssumePrime = 1;
	end	else if (num==16'd56081) begin
		AssumePrime = 1;
	end	else if (num==16'd56087) begin
		AssumePrime = 1;
	end	else if (num==16'd56093) begin
		AssumePrime = 1;
	end	else if (num==16'd56099) begin
		AssumePrime = 1;
	end	else if (num==16'd56101) begin
		AssumePrime = 1;
	end	else if (num==16'd56113) begin
		AssumePrime = 1;
	end	else if (num==16'd56123) begin
		AssumePrime = 1;
	end	else if (num==16'd56131) begin
		AssumePrime = 1;
	end	else if (num==16'd56149) begin
		AssumePrime = 1;
	end	else if (num==16'd56167) begin
		AssumePrime = 1;
	end	else if (num==16'd56171) begin
		AssumePrime = 1;
	end	else if (num==16'd56179) begin
		AssumePrime = 1;
	end	else if (num==16'd56197) begin
		AssumePrime = 1;
	end	else if (num==16'd56207) begin
		AssumePrime = 1;
	end	else if (num==16'd56209) begin
		AssumePrime = 1;
	end	else if (num==16'd56237) begin
		AssumePrime = 1;
	end	else if (num==16'd56239) begin
		AssumePrime = 1;
	end	else if (num==16'd56249) begin
		AssumePrime = 1;
	end	else if (num==16'd56263) begin
		AssumePrime = 1;
	end	else if (num==16'd56267) begin
		AssumePrime = 1;
	end	else if (num==16'd56269) begin
		AssumePrime = 1;
	end	else if (num==16'd56299) begin
		AssumePrime = 1;
	end	else if (num==16'd56311) begin
		AssumePrime = 1;
	end	else if (num==16'd56333) begin
		AssumePrime = 1;
	end	else if (num==16'd56359) begin
		AssumePrime = 1;
	end	else if (num==16'd56369) begin
		AssumePrime = 1;
	end	else if (num==16'd56377) begin
		AssumePrime = 1;
	end	else if (num==16'd56383) begin
		AssumePrime = 1;
	end	else if (num==16'd56393) begin
		AssumePrime = 1;
	end	else if (num==16'd56401) begin
		AssumePrime = 1;
	end	else if (num==16'd56417) begin
		AssumePrime = 1;
	end	else if (num==16'd56431) begin
		AssumePrime = 1;
	end	else if (num==16'd56437) begin
		AssumePrime = 1;
	end	else if (num==16'd56443) begin
		AssumePrime = 1;
	end	else if (num==16'd56453) begin
		AssumePrime = 1;
	end	else if (num==16'd56467) begin
		AssumePrime = 1;
	end	else if (num==16'd56473) begin
		AssumePrime = 1;
	end	else if (num==16'd56477) begin
		AssumePrime = 1;
	end	else if (num==16'd56479) begin
		AssumePrime = 1;
	end	else if (num==16'd56489) begin
		AssumePrime = 1;
	end	else if (num==16'd56501) begin
		AssumePrime = 1;
	end	else if (num==16'd56503) begin
		AssumePrime = 1;
	end	else if (num==16'd56509) begin
		AssumePrime = 1;
	end	else if (num==16'd56519) begin
		AssumePrime = 1;
	end	else if (num==16'd56527) begin
		AssumePrime = 1;
	end	else if (num==16'd56531) begin
		AssumePrime = 1;
	end	else if (num==16'd56533) begin
		AssumePrime = 1;
	end	else if (num==16'd56543) begin
		AssumePrime = 1;
	end	else if (num==16'd56569) begin
		AssumePrime = 1;
	end	else if (num==16'd56591) begin
		AssumePrime = 1;
	end	else if (num==16'd56597) begin
		AssumePrime = 1;
	end	else if (num==16'd56599) begin
		AssumePrime = 1;
	end	else if (num==16'd56611) begin
		AssumePrime = 1;
	end	else if (num==16'd56629) begin
		AssumePrime = 1;
	end	else if (num==16'd56633) begin
		AssumePrime = 1;
	end	else if (num==16'd56659) begin
		AssumePrime = 1;
	end	else if (num==16'd56663) begin
		AssumePrime = 1;
	end	else if (num==16'd56671) begin
		AssumePrime = 1;
	end	else if (num==16'd56681) begin
		AssumePrime = 1;
	end	else if (num==16'd56687) begin
		AssumePrime = 1;
	end	else if (num==16'd56701) begin
		AssumePrime = 1;
	end	else if (num==16'd56711) begin
		AssumePrime = 1;
	end	else if (num==16'd56713) begin
		AssumePrime = 1;
	end	else if (num==16'd56731) begin
		AssumePrime = 1;
	end	else if (num==16'd56737) begin
		AssumePrime = 1;
	end	else if (num==16'd56747) begin
		AssumePrime = 1;
	end	else if (num==16'd56767) begin
		AssumePrime = 1;
	end	else if (num==16'd56773) begin
		AssumePrime = 1;
	end	else if (num==16'd56779) begin
		AssumePrime = 1;
	end	else if (num==16'd56783) begin
		AssumePrime = 1;
	end	else if (num==16'd56807) begin
		AssumePrime = 1;
	end	else if (num==16'd56809) begin
		AssumePrime = 1;
	end	else if (num==16'd56813) begin
		AssumePrime = 1;
	end	else if (num==16'd56821) begin
		AssumePrime = 1;
	end	else if (num==16'd56827) begin
		AssumePrime = 1;
	end	else if (num==16'd56843) begin
		AssumePrime = 1;
	end	else if (num==16'd56857) begin
		AssumePrime = 1;
	end	else if (num==16'd56873) begin
		AssumePrime = 1;
	end	else if (num==16'd56891) begin
		AssumePrime = 1;
	end	else if (num==16'd56893) begin
		AssumePrime = 1;
	end	else if (num==16'd56897) begin
		AssumePrime = 1;
	end	else if (num==16'd56909) begin
		AssumePrime = 1;
	end	else if (num==16'd56911) begin
		AssumePrime = 1;
	end	else if (num==16'd56921) begin
		AssumePrime = 1;
	end	else if (num==16'd56923) begin
		AssumePrime = 1;
	end	else if (num==16'd56929) begin
		AssumePrime = 1;
	end	else if (num==16'd56941) begin
		AssumePrime = 1;
	end	else if (num==16'd56951) begin
		AssumePrime = 1;
	end	else if (num==16'd56957) begin
		AssumePrime = 1;
	end	else if (num==16'd56963) begin
		AssumePrime = 1;
	end	else if (num==16'd56983) begin
		AssumePrime = 1;
	end	else if (num==16'd56989) begin
		AssumePrime = 1;
	end	else if (num==16'd56993) begin
		AssumePrime = 1;
	end	else if (num==16'd56999) begin
		AssumePrime = 1;
	end	else if (num==16'd57037) begin
		AssumePrime = 1;
	end	else if (num==16'd57041) begin
		AssumePrime = 1;
	end	else if (num==16'd57047) begin
		AssumePrime = 1;
	end	else if (num==16'd57059) begin
		AssumePrime = 1;
	end	else if (num==16'd57073) begin
		AssumePrime = 1;
	end	else if (num==16'd57077) begin
		AssumePrime = 1;
	end	else if (num==16'd57089) begin
		AssumePrime = 1;
	end	else if (num==16'd57097) begin
		AssumePrime = 1;
	end	else if (num==16'd57107) begin
		AssumePrime = 1;
	end	else if (num==16'd57119) begin
		AssumePrime = 1;
	end	else if (num==16'd57131) begin
		AssumePrime = 1;
	end	else if (num==16'd57139) begin
		AssumePrime = 1;
	end	else if (num==16'd57143) begin
		AssumePrime = 1;
	end	else if (num==16'd57149) begin
		AssumePrime = 1;
	end	else if (num==16'd57163) begin
		AssumePrime = 1;
	end	else if (num==16'd57173) begin
		AssumePrime = 1;
	end	else if (num==16'd57179) begin
		AssumePrime = 1;
	end	else if (num==16'd57191) begin
		AssumePrime = 1;
	end	else if (num==16'd57193) begin
		AssumePrime = 1;
	end	else if (num==16'd57203) begin
		AssumePrime = 1;
	end	else if (num==16'd57221) begin
		AssumePrime = 1;
	end	else if (num==16'd57223) begin
		AssumePrime = 1;
	end	else if (num==16'd57241) begin
		AssumePrime = 1;
	end	else if (num==16'd57251) begin
		AssumePrime = 1;
	end	else if (num==16'd57259) begin
		AssumePrime = 1;
	end	else if (num==16'd57269) begin
		AssumePrime = 1;
	end	else if (num==16'd57271) begin
		AssumePrime = 1;
	end	else if (num==16'd57283) begin
		AssumePrime = 1;
	end	else if (num==16'd57287) begin
		AssumePrime = 1;
	end	else if (num==16'd57301) begin
		AssumePrime = 1;
	end	else if (num==16'd57329) begin
		AssumePrime = 1;
	end	else if (num==16'd57331) begin
		AssumePrime = 1;
	end	else if (num==16'd57347) begin
		AssumePrime = 1;
	end	else if (num==16'd57349) begin
		AssumePrime = 1;
	end	else if (num==16'd57367) begin
		AssumePrime = 1;
	end	else if (num==16'd57373) begin
		AssumePrime = 1;
	end	else if (num==16'd57383) begin
		AssumePrime = 1;
	end	else if (num==16'd57389) begin
		AssumePrime = 1;
	end	else if (num==16'd57397) begin
		AssumePrime = 1;
	end	else if (num==16'd57413) begin
		AssumePrime = 1;
	end	else if (num==16'd57427) begin
		AssumePrime = 1;
	end	else if (num==16'd57457) begin
		AssumePrime = 1;
	end	else if (num==16'd57467) begin
		AssumePrime = 1;
	end	else if (num==16'd57487) begin
		AssumePrime = 1;
	end	else if (num==16'd57493) begin
		AssumePrime = 1;
	end	else if (num==16'd57503) begin
		AssumePrime = 1;
	end	else if (num==16'd57527) begin
		AssumePrime = 1;
	end	else if (num==16'd57529) begin
		AssumePrime = 1;
	end	else if (num==16'd57557) begin
		AssumePrime = 1;
	end	else if (num==16'd57559) begin
		AssumePrime = 1;
	end	else if (num==16'd57571) begin
		AssumePrime = 1;
	end	else if (num==16'd57587) begin
		AssumePrime = 1;
	end	else if (num==16'd57593) begin
		AssumePrime = 1;
	end	else if (num==16'd57601) begin
		AssumePrime = 1;
	end	else if (num==16'd57637) begin
		AssumePrime = 1;
	end	else if (num==16'd57641) begin
		AssumePrime = 1;
	end	else if (num==16'd57649) begin
		AssumePrime = 1;
	end	else if (num==16'd57653) begin
		AssumePrime = 1;
	end	else if (num==16'd57667) begin
		AssumePrime = 1;
	end	else if (num==16'd57679) begin
		AssumePrime = 1;
	end	else if (num==16'd57689) begin
		AssumePrime = 1;
	end	else if (num==16'd57697) begin
		AssumePrime = 1;
	end	else if (num==16'd57709) begin
		AssumePrime = 1;
	end	else if (num==16'd57713) begin
		AssumePrime = 1;
	end	else if (num==16'd57719) begin
		AssumePrime = 1;
	end	else if (num==16'd57727) begin
		AssumePrime = 1;
	end	else if (num==16'd57731) begin
		AssumePrime = 1;
	end	else if (num==16'd57737) begin
		AssumePrime = 1;
	end	else if (num==16'd57751) begin
		AssumePrime = 1;
	end	else if (num==16'd57773) begin
		AssumePrime = 1;
	end	else if (num==16'd57781) begin
		AssumePrime = 1;
	end	else if (num==16'd57787) begin
		AssumePrime = 1;
	end	else if (num==16'd57791) begin
		AssumePrime = 1;
	end	else if (num==16'd57793) begin
		AssumePrime = 1;
	end	else if (num==16'd57803) begin
		AssumePrime = 1;
	end	else if (num==16'd57809) begin
		AssumePrime = 1;
	end	else if (num==16'd57829) begin
		AssumePrime = 1;
	end	else if (num==16'd57839) begin
		AssumePrime = 1;
	end	else if (num==16'd57847) begin
		AssumePrime = 1;
	end	else if (num==16'd57853) begin
		AssumePrime = 1;
	end	else if (num==16'd57859) begin
		AssumePrime = 1;
	end	else if (num==16'd57881) begin
		AssumePrime = 1;
	end	else if (num==16'd57899) begin
		AssumePrime = 1;
	end	else if (num==16'd57901) begin
		AssumePrime = 1;
	end	else if (num==16'd57917) begin
		AssumePrime = 1;
	end	else if (num==16'd57923) begin
		AssumePrime = 1;
	end	else if (num==16'd57943) begin
		AssumePrime = 1;
	end	else if (num==16'd57947) begin
		AssumePrime = 1;
	end	else if (num==16'd57973) begin
		AssumePrime = 1;
	end	else if (num==16'd57977) begin
		AssumePrime = 1;
	end	else if (num==16'd57991) begin
		AssumePrime = 1;
	end	else if (num==16'd58013) begin
		AssumePrime = 1;
	end	else if (num==16'd58027) begin
		AssumePrime = 1;
	end	else if (num==16'd58031) begin
		AssumePrime = 1;
	end	else if (num==16'd58043) begin
		AssumePrime = 1;
	end	else if (num==16'd58049) begin
		AssumePrime = 1;
	end	else if (num==16'd58057) begin
		AssumePrime = 1;
	end	else if (num==16'd58061) begin
		AssumePrime = 1;
	end	else if (num==16'd58067) begin
		AssumePrime = 1;
	end	else if (num==16'd58073) begin
		AssumePrime = 1;
	end	else if (num==16'd58099) begin
		AssumePrime = 1;
	end	else if (num==16'd58109) begin
		AssumePrime = 1;
	end	else if (num==16'd58111) begin
		AssumePrime = 1;
	end	else if (num==16'd58129) begin
		AssumePrime = 1;
	end	else if (num==16'd58147) begin
		AssumePrime = 1;
	end	else if (num==16'd58151) begin
		AssumePrime = 1;
	end	else if (num==16'd58153) begin
		AssumePrime = 1;
	end	else if (num==16'd58169) begin
		AssumePrime = 1;
	end	else if (num==16'd58171) begin
		AssumePrime = 1;
	end	else if (num==16'd58189) begin
		AssumePrime = 1;
	end	else if (num==16'd58193) begin
		AssumePrime = 1;
	end	else if (num==16'd58199) begin
		AssumePrime = 1;
	end	else if (num==16'd58207) begin
		AssumePrime = 1;
	end	else if (num==16'd58211) begin
		AssumePrime = 1;
	end	else if (num==16'd58217) begin
		AssumePrime = 1;
	end	else if (num==16'd58229) begin
		AssumePrime = 1;
	end	else if (num==16'd58231) begin
		AssumePrime = 1;
	end	else if (num==16'd58237) begin
		AssumePrime = 1;
	end	else if (num==16'd58243) begin
		AssumePrime = 1;
	end	else if (num==16'd58271) begin
		AssumePrime = 1;
	end	else if (num==16'd58309) begin
		AssumePrime = 1;
	end	else if (num==16'd58313) begin
		AssumePrime = 1;
	end	else if (num==16'd58321) begin
		AssumePrime = 1;
	end	else if (num==16'd58337) begin
		AssumePrime = 1;
	end	else if (num==16'd58363) begin
		AssumePrime = 1;
	end	else if (num==16'd58367) begin
		AssumePrime = 1;
	end	else if (num==16'd58369) begin
		AssumePrime = 1;
	end	else if (num==16'd58379) begin
		AssumePrime = 1;
	end	else if (num==16'd58391) begin
		AssumePrime = 1;
	end	else if (num==16'd58393) begin
		AssumePrime = 1;
	end	else if (num==16'd58403) begin
		AssumePrime = 1;
	end	else if (num==16'd58411) begin
		AssumePrime = 1;
	end	else if (num==16'd58417) begin
		AssumePrime = 1;
	end	else if (num==16'd58427) begin
		AssumePrime = 1;
	end	else if (num==16'd58439) begin
		AssumePrime = 1;
	end	else if (num==16'd58441) begin
		AssumePrime = 1;
	end	else if (num==16'd58451) begin
		AssumePrime = 1;
	end	else if (num==16'd58453) begin
		AssumePrime = 1;
	end	else if (num==16'd58477) begin
		AssumePrime = 1;
	end	else if (num==16'd58481) begin
		AssumePrime = 1;
	end	else if (num==16'd58511) begin
		AssumePrime = 1;
	end	else if (num==16'd58537) begin
		AssumePrime = 1;
	end	else if (num==16'd58543) begin
		AssumePrime = 1;
	end	else if (num==16'd58549) begin
		AssumePrime = 1;
	end	else if (num==16'd58567) begin
		AssumePrime = 1;
	end	else if (num==16'd58573) begin
		AssumePrime = 1;
	end	else if (num==16'd58579) begin
		AssumePrime = 1;
	end	else if (num==16'd58601) begin
		AssumePrime = 1;
	end	else if (num==16'd58603) begin
		AssumePrime = 1;
	end	else if (num==16'd58613) begin
		AssumePrime = 1;
	end	else if (num==16'd58631) begin
		AssumePrime = 1;
	end	else if (num==16'd58657) begin
		AssumePrime = 1;
	end	else if (num==16'd58661) begin
		AssumePrime = 1;
	end	else if (num==16'd58679) begin
		AssumePrime = 1;
	end	else if (num==16'd58687) begin
		AssumePrime = 1;
	end	else if (num==16'd58693) begin
		AssumePrime = 1;
	end	else if (num==16'd58699) begin
		AssumePrime = 1;
	end	else if (num==16'd58711) begin
		AssumePrime = 1;
	end	else if (num==16'd58727) begin
		AssumePrime = 1;
	end	else if (num==16'd58733) begin
		AssumePrime = 1;
	end	else if (num==16'd58741) begin
		AssumePrime = 1;
	end	else if (num==16'd58757) begin
		AssumePrime = 1;
	end	else if (num==16'd58763) begin
		AssumePrime = 1;
	end	else if (num==16'd58771) begin
		AssumePrime = 1;
	end	else if (num==16'd58787) begin
		AssumePrime = 1;
	end	else if (num==16'd58789) begin
		AssumePrime = 1;
	end	else if (num==16'd58831) begin
		AssumePrime = 1;
	end	else if (num==16'd58889) begin
		AssumePrime = 1;
	end	else if (num==16'd58897) begin
		AssumePrime = 1;
	end	else if (num==16'd58901) begin
		AssumePrime = 1;
	end	else if (num==16'd58907) begin
		AssumePrime = 1;
	end	else if (num==16'd58909) begin
		AssumePrime = 1;
	end	else if (num==16'd58913) begin
		AssumePrime = 1;
	end	else if (num==16'd58921) begin
		AssumePrime = 1;
	end	else if (num==16'd58937) begin
		AssumePrime = 1;
	end	else if (num==16'd58943) begin
		AssumePrime = 1;
	end	else if (num==16'd58963) begin
		AssumePrime = 1;
	end	else if (num==16'd58967) begin
		AssumePrime = 1;
	end	else if (num==16'd58979) begin
		AssumePrime = 1;
	end	else if (num==16'd58991) begin
		AssumePrime = 1;
	end	else if (num==16'd58997) begin
		AssumePrime = 1;
	end	else if (num==16'd59009) begin
		AssumePrime = 1;
	end	else if (num==16'd59011) begin
		AssumePrime = 1;
	end	else if (num==16'd59021) begin
		AssumePrime = 1;
	end	else if (num==16'd59023) begin
		AssumePrime = 1;
	end	else if (num==16'd59029) begin
		AssumePrime = 1;
	end	else if (num==16'd59051) begin
		AssumePrime = 1;
	end	else if (num==16'd59053) begin
		AssumePrime = 1;
	end	else if (num==16'd59063) begin
		AssumePrime = 1;
	end	else if (num==16'd59069) begin
		AssumePrime = 1;
	end	else if (num==16'd59077) begin
		AssumePrime = 1;
	end	else if (num==16'd59083) begin
		AssumePrime = 1;
	end	else if (num==16'd59093) begin
		AssumePrime = 1;
	end	else if (num==16'd59107) begin
		AssumePrime = 1;
	end	else if (num==16'd59113) begin
		AssumePrime = 1;
	end	else if (num==16'd59119) begin
		AssumePrime = 1;
	end	else if (num==16'd59123) begin
		AssumePrime = 1;
	end	else if (num==16'd59141) begin
		AssumePrime = 1;
	end	else if (num==16'd59149) begin
		AssumePrime = 1;
	end	else if (num==16'd59159) begin
		AssumePrime = 1;
	end	else if (num==16'd59167) begin
		AssumePrime = 1;
	end	else if (num==16'd59183) begin
		AssumePrime = 1;
	end	else if (num==16'd59197) begin
		AssumePrime = 1;
	end	else if (num==16'd59207) begin
		AssumePrime = 1;
	end	else if (num==16'd59209) begin
		AssumePrime = 1;
	end	else if (num==16'd59219) begin
		AssumePrime = 1;
	end	else if (num==16'd59221) begin
		AssumePrime = 1;
	end	else if (num==16'd59233) begin
		AssumePrime = 1;
	end	else if (num==16'd59239) begin
		AssumePrime = 1;
	end	else if (num==16'd59243) begin
		AssumePrime = 1;
	end	else if (num==16'd59263) begin
		AssumePrime = 1;
	end	else if (num==16'd59273) begin
		AssumePrime = 1;
	end	else if (num==16'd59281) begin
		AssumePrime = 1;
	end	else if (num==16'd59333) begin
		AssumePrime = 1;
	end	else if (num==16'd59341) begin
		AssumePrime = 1;
	end	else if (num==16'd59351) begin
		AssumePrime = 1;
	end	else if (num==16'd59357) begin
		AssumePrime = 1;
	end	else if (num==16'd59359) begin
		AssumePrime = 1;
	end	else if (num==16'd59369) begin
		AssumePrime = 1;
	end	else if (num==16'd59377) begin
		AssumePrime = 1;
	end	else if (num==16'd59387) begin
		AssumePrime = 1;
	end	else if (num==16'd59393) begin
		AssumePrime = 1;
	end	else if (num==16'd59399) begin
		AssumePrime = 1;
	end	else if (num==16'd59407) begin
		AssumePrime = 1;
	end	else if (num==16'd59417) begin
		AssumePrime = 1;
	end	else if (num==16'd59419) begin
		AssumePrime = 1;
	end	else if (num==16'd59441) begin
		AssumePrime = 1;
	end	else if (num==16'd59443) begin
		AssumePrime = 1;
	end	else if (num==16'd59447) begin
		AssumePrime = 1;
	end	else if (num==16'd59453) begin
		AssumePrime = 1;
	end	else if (num==16'd59467) begin
		AssumePrime = 1;
	end	else if (num==16'd59471) begin
		AssumePrime = 1;
	end	else if (num==16'd59473) begin
		AssumePrime = 1;
	end	else if (num==16'd59497) begin
		AssumePrime = 1;
	end	else if (num==16'd59509) begin
		AssumePrime = 1;
	end	else if (num==16'd59513) begin
		AssumePrime = 1;
	end	else if (num==16'd59539) begin
		AssumePrime = 1;
	end	else if (num==16'd59557) begin
		AssumePrime = 1;
	end	else if (num==16'd59561) begin
		AssumePrime = 1;
	end	else if (num==16'd59567) begin
		AssumePrime = 1;
	end	else if (num==16'd59581) begin
		AssumePrime = 1;
	end	else if (num==16'd59611) begin
		AssumePrime = 1;
	end	else if (num==16'd59617) begin
		AssumePrime = 1;
	end	else if (num==16'd59621) begin
		AssumePrime = 1;
	end	else if (num==16'd59627) begin
		AssumePrime = 1;
	end	else if (num==16'd59629) begin
		AssumePrime = 1;
	end	else if (num==16'd59651) begin
		AssumePrime = 1;
	end	else if (num==16'd59659) begin
		AssumePrime = 1;
	end	else if (num==16'd59663) begin
		AssumePrime = 1;
	end	else if (num==16'd59669) begin
		AssumePrime = 1;
	end	else if (num==16'd59671) begin
		AssumePrime = 1;
	end	else if (num==16'd59693) begin
		AssumePrime = 1;
	end	else if (num==16'd59699) begin
		AssumePrime = 1;
	end	else if (num==16'd59707) begin
		AssumePrime = 1;
	end	else if (num==16'd59723) begin
		AssumePrime = 1;
	end	else if (num==16'd59729) begin
		AssumePrime = 1;
	end	else if (num==16'd59743) begin
		AssumePrime = 1;
	end	else if (num==16'd59747) begin
		AssumePrime = 1;
	end	else if (num==16'd59753) begin
		AssumePrime = 1;
	end	else if (num==16'd59771) begin
		AssumePrime = 1;
	end	else if (num==16'd59779) begin
		AssumePrime = 1;
	end	else if (num==16'd59791) begin
		AssumePrime = 1;
	end	else if (num==16'd59797) begin
		AssumePrime = 1;
	end	else if (num==16'd59809) begin
		AssumePrime = 1;
	end	else if (num==16'd59833) begin
		AssumePrime = 1;
	end	else if (num==16'd59863) begin
		AssumePrime = 1;
	end	else if (num==16'd59879) begin
		AssumePrime = 1;
	end	else if (num==16'd59887) begin
		AssumePrime = 1;
	end	else if (num==16'd59921) begin
		AssumePrime = 1;
	end	else if (num==16'd59929) begin
		AssumePrime = 1;
	end	else if (num==16'd59951) begin
		AssumePrime = 1;
	end	else if (num==16'd59957) begin
		AssumePrime = 1;
	end	else if (num==16'd59971) begin
		AssumePrime = 1;
	end	else if (num==16'd59981) begin
		AssumePrime = 1;
	end	else if (num==16'd59999) begin
		AssumePrime = 1;
	end	else if (num==16'd60013) begin
		AssumePrime = 1;
	end	else if (num==16'd60017) begin
		AssumePrime = 1;
	end	else if (num==16'd60029) begin
		AssumePrime = 1;
	end	else if (num==16'd60037) begin
		AssumePrime = 1;
	end	else if (num==16'd60041) begin
		AssumePrime = 1;
	end	else if (num==16'd60077) begin
		AssumePrime = 1;
	end	else if (num==16'd60083) begin
		AssumePrime = 1;
	end	else if (num==16'd60089) begin
		AssumePrime = 1;
	end	else if (num==16'd60091) begin
		AssumePrime = 1;
	end	else if (num==16'd60101) begin
		AssumePrime = 1;
	end	else if (num==16'd60103) begin
		AssumePrime = 1;
	end	else if (num==16'd60107) begin
		AssumePrime = 1;
	end	else if (num==16'd60127) begin
		AssumePrime = 1;
	end	else if (num==16'd60133) begin
		AssumePrime = 1;
	end	else if (num==16'd60139) begin
		AssumePrime = 1;
	end	else if (num==16'd60149) begin
		AssumePrime = 1;
	end	else if (num==16'd60161) begin
		AssumePrime = 1;
	end	else if (num==16'd60167) begin
		AssumePrime = 1;
	end	else if (num==16'd60169) begin
		AssumePrime = 1;
	end	else if (num==16'd60209) begin
		AssumePrime = 1;
	end	else if (num==16'd60217) begin
		AssumePrime = 1;
	end	else if (num==16'd60223) begin
		AssumePrime = 1;
	end	else if (num==16'd60251) begin
		AssumePrime = 1;
	end	else if (num==16'd60257) begin
		AssumePrime = 1;
	end	else if (num==16'd60259) begin
		AssumePrime = 1;
	end	else if (num==16'd60271) begin
		AssumePrime = 1;
	end	else if (num==16'd60289) begin
		AssumePrime = 1;
	end	else if (num==16'd60293) begin
		AssumePrime = 1;
	end	else if (num==16'd60317) begin
		AssumePrime = 1;
	end	else if (num==16'd60331) begin
		AssumePrime = 1;
	end	else if (num==16'd60337) begin
		AssumePrime = 1;
	end	else if (num==16'd60343) begin
		AssumePrime = 1;
	end	else if (num==16'd60353) begin
		AssumePrime = 1;
	end	else if (num==16'd60373) begin
		AssumePrime = 1;
	end	else if (num==16'd60383) begin
		AssumePrime = 1;
	end	else if (num==16'd60397) begin
		AssumePrime = 1;
	end	else if (num==16'd60413) begin
		AssumePrime = 1;
	end	else if (num==16'd60427) begin
		AssumePrime = 1;
	end	else if (num==16'd60443) begin
		AssumePrime = 1;
	end	else if (num==16'd60449) begin
		AssumePrime = 1;
	end	else if (num==16'd60457) begin
		AssumePrime = 1;
	end	else if (num==16'd60493) begin
		AssumePrime = 1;
	end	else if (num==16'd60497) begin
		AssumePrime = 1;
	end	else if (num==16'd60509) begin
		AssumePrime = 1;
	end	else if (num==16'd60521) begin
		AssumePrime = 1;
	end	else if (num==16'd60527) begin
		AssumePrime = 1;
	end	else if (num==16'd60539) begin
		AssumePrime = 1;
	end	else if (num==16'd60589) begin
		AssumePrime = 1;
	end	else if (num==16'd60601) begin
		AssumePrime = 1;
	end	else if (num==16'd60607) begin
		AssumePrime = 1;
	end	else if (num==16'd60611) begin
		AssumePrime = 1;
	end	else if (num==16'd60617) begin
		AssumePrime = 1;
	end	else if (num==16'd60623) begin
		AssumePrime = 1;
	end	else if (num==16'd60631) begin
		AssumePrime = 1;
	end	else if (num==16'd60637) begin
		AssumePrime = 1;
	end	else if (num==16'd60647) begin
		AssumePrime = 1;
	end	else if (num==16'd60649) begin
		AssumePrime = 1;
	end	else if (num==16'd60659) begin
		AssumePrime = 1;
	end	else if (num==16'd60661) begin
		AssumePrime = 1;
	end	else if (num==16'd60679) begin
		AssumePrime = 1;
	end	else if (num==16'd60689) begin
		AssumePrime = 1;
	end	else if (num==16'd60703) begin
		AssumePrime = 1;
	end	else if (num==16'd60719) begin
		AssumePrime = 1;
	end	else if (num==16'd60727) begin
		AssumePrime = 1;
	end	else if (num==16'd60733) begin
		AssumePrime = 1;
	end	else if (num==16'd60737) begin
		AssumePrime = 1;
	end	else if (num==16'd60757) begin
		AssumePrime = 1;
	end	else if (num==16'd60761) begin
		AssumePrime = 1;
	end	else if (num==16'd60763) begin
		AssumePrime = 1;
	end	else if (num==16'd60773) begin
		AssumePrime = 1;
	end	else if (num==16'd60779) begin
		AssumePrime = 1;
	end	else if (num==16'd60793) begin
		AssumePrime = 1;
	end	else if (num==16'd60811) begin
		AssumePrime = 1;
	end	else if (num==16'd60821) begin
		AssumePrime = 1;
	end	else if (num==16'd60859) begin
		AssumePrime = 1;
	end	else if (num==16'd60869) begin
		AssumePrime = 1;
	end	else if (num==16'd60887) begin
		AssumePrime = 1;
	end	else if (num==16'd60889) begin
		AssumePrime = 1;
	end	else if (num==16'd60899) begin
		AssumePrime = 1;
	end	else if (num==16'd60901) begin
		AssumePrime = 1;
	end	else if (num==16'd60913) begin
		AssumePrime = 1;
	end	else if (num==16'd60917) begin
		AssumePrime = 1;
	end	else if (num==16'd60919) begin
		AssumePrime = 1;
	end	else if (num==16'd60923) begin
		AssumePrime = 1;
	end	else if (num==16'd60937) begin
		AssumePrime = 1;
	end	else if (num==16'd60943) begin
		AssumePrime = 1;
	end	else if (num==16'd60953) begin
		AssumePrime = 1;
	end	else if (num==16'd60961) begin
		AssumePrime = 1;
	end	else if (num==16'd61001) begin
		AssumePrime = 1;
	end	else if (num==16'd61007) begin
		AssumePrime = 1;
	end	else if (num==16'd61027) begin
		AssumePrime = 1;
	end	else if (num==16'd61031) begin
		AssumePrime = 1;
	end	else if (num==16'd61043) begin
		AssumePrime = 1;
	end	else if (num==16'd61051) begin
		AssumePrime = 1;
	end	else if (num==16'd61057) begin
		AssumePrime = 1;
	end	else if (num==16'd61091) begin
		AssumePrime = 1;
	end	else if (num==16'd61099) begin
		AssumePrime = 1;
	end	else if (num==16'd61121) begin
		AssumePrime = 1;
	end	else if (num==16'd61129) begin
		AssumePrime = 1;
	end	else if (num==16'd61141) begin
		AssumePrime = 1;
	end	else if (num==16'd61151) begin
		AssumePrime = 1;
	end	else if (num==16'd61153) begin
		AssumePrime = 1;
	end	else if (num==16'd61169) begin
		AssumePrime = 1;
	end	else if (num==16'd61211) begin
		AssumePrime = 1;
	end	else if (num==16'd61223) begin
		AssumePrime = 1;
	end	else if (num==16'd61231) begin
		AssumePrime = 1;
	end	else if (num==16'd61253) begin
		AssumePrime = 1;
	end	else if (num==16'd61261) begin
		AssumePrime = 1;
	end	else if (num==16'd61283) begin
		AssumePrime = 1;
	end	else if (num==16'd61291) begin
		AssumePrime = 1;
	end	else if (num==16'd61297) begin
		AssumePrime = 1;
	end	else if (num==16'd61331) begin
		AssumePrime = 1;
	end	else if (num==16'd61333) begin
		AssumePrime = 1;
	end	else if (num==16'd61339) begin
		AssumePrime = 1;
	end	else if (num==16'd61343) begin
		AssumePrime = 1;
	end	else if (num==16'd61357) begin
		AssumePrime = 1;
	end	else if (num==16'd61363) begin
		AssumePrime = 1;
	end	else if (num==16'd61379) begin
		AssumePrime = 1;
	end	else if (num==16'd61381) begin
		AssumePrime = 1;
	end	else if (num==16'd61403) begin
		AssumePrime = 1;
	end	else if (num==16'd61409) begin
		AssumePrime = 1;
	end	else if (num==16'd61417) begin
		AssumePrime = 1;
	end	else if (num==16'd61441) begin
		AssumePrime = 1;
	end	else if (num==16'd61463) begin
		AssumePrime = 1;
	end	else if (num==16'd61469) begin
		AssumePrime = 1;
	end	else if (num==16'd61471) begin
		AssumePrime = 1;
	end	else if (num==16'd61483) begin
		AssumePrime = 1;
	end	else if (num==16'd61487) begin
		AssumePrime = 1;
	end	else if (num==16'd61493) begin
		AssumePrime = 1;
	end	else if (num==16'd61507) begin
		AssumePrime = 1;
	end	else if (num==16'd61511) begin
		AssumePrime = 1;
	end	else if (num==16'd61519) begin
		AssumePrime = 1;
	end	else if (num==16'd61543) begin
		AssumePrime = 1;
	end	else if (num==16'd61547) begin
		AssumePrime = 1;
	end	else if (num==16'd61553) begin
		AssumePrime = 1;
	end	else if (num==16'd61559) begin
		AssumePrime = 1;
	end	else if (num==16'd61561) begin
		AssumePrime = 1;
	end	else if (num==16'd61583) begin
		AssumePrime = 1;
	end	else if (num==16'd61603) begin
		AssumePrime = 1;
	end	else if (num==16'd61609) begin
		AssumePrime = 1;
	end	else if (num==16'd61613) begin
		AssumePrime = 1;
	end	else if (num==16'd61627) begin
		AssumePrime = 1;
	end	else if (num==16'd61631) begin
		AssumePrime = 1;
	end	else if (num==16'd61637) begin
		AssumePrime = 1;
	end	else if (num==16'd61643) begin
		AssumePrime = 1;
	end	else if (num==16'd61651) begin
		AssumePrime = 1;
	end	else if (num==16'd61657) begin
		AssumePrime = 1;
	end	else if (num==16'd61667) begin
		AssumePrime = 1;
	end	else if (num==16'd61673) begin
		AssumePrime = 1;
	end	else if (num==16'd61681) begin
		AssumePrime = 1;
	end	else if (num==16'd61687) begin
		AssumePrime = 1;
	end	else if (num==16'd61703) begin
		AssumePrime = 1;
	end	else if (num==16'd61717) begin
		AssumePrime = 1;
	end	else if (num==16'd61723) begin
		AssumePrime = 1;
	end	else if (num==16'd61729) begin
		AssumePrime = 1;
	end	else if (num==16'd61751) begin
		AssumePrime = 1;
	end	else if (num==16'd61757) begin
		AssumePrime = 1;
	end	else if (num==16'd61781) begin
		AssumePrime = 1;
	end	else if (num==16'd61813) begin
		AssumePrime = 1;
	end	else if (num==16'd61819) begin
		AssumePrime = 1;
	end	else if (num==16'd61837) begin
		AssumePrime = 1;
	end	else if (num==16'd61843) begin
		AssumePrime = 1;
	end	else if (num==16'd61861) begin
		AssumePrime = 1;
	end	else if (num==16'd61871) begin
		AssumePrime = 1;
	end	else if (num==16'd61879) begin
		AssumePrime = 1;
	end	else if (num==16'd61909) begin
		AssumePrime = 1;
	end	else if (num==16'd61927) begin
		AssumePrime = 1;
	end	else if (num==16'd61933) begin
		AssumePrime = 1;
	end	else if (num==16'd61949) begin
		AssumePrime = 1;
	end	else if (num==16'd61961) begin
		AssumePrime = 1;
	end	else if (num==16'd61967) begin
		AssumePrime = 1;
	end	else if (num==16'd61979) begin
		AssumePrime = 1;
	end	else if (num==16'd61981) begin
		AssumePrime = 1;
	end	else if (num==16'd61987) begin
		AssumePrime = 1;
	end	else if (num==16'd61991) begin
		AssumePrime = 1;
	end	else if (num==16'd62003) begin
		AssumePrime = 1;
	end	else if (num==16'd62011) begin
		AssumePrime = 1;
	end	else if (num==16'd62017) begin
		AssumePrime = 1;
	end	else if (num==16'd62039) begin
		AssumePrime = 1;
	end	else if (num==16'd62047) begin
		AssumePrime = 1;
	end	else if (num==16'd62053) begin
		AssumePrime = 1;
	end	else if (num==16'd62057) begin
		AssumePrime = 1;
	end	else if (num==16'd62071) begin
		AssumePrime = 1;
	end	else if (num==16'd62081) begin
		AssumePrime = 1;
	end	else if (num==16'd62099) begin
		AssumePrime = 1;
	end	else if (num==16'd62119) begin
		AssumePrime = 1;
	end	else if (num==16'd62129) begin
		AssumePrime = 1;
	end	else if (num==16'd62131) begin
		AssumePrime = 1;
	end	else if (num==16'd62137) begin
		AssumePrime = 1;
	end	else if (num==16'd62141) begin
		AssumePrime = 1;
	end	else if (num==16'd62143) begin
		AssumePrime = 1;
	end	else if (num==16'd62171) begin
		AssumePrime = 1;
	end	else if (num==16'd62189) begin
		AssumePrime = 1;
	end	else if (num==16'd62191) begin
		AssumePrime = 1;
	end	else if (num==16'd62201) begin
		AssumePrime = 1;
	end	else if (num==16'd62207) begin
		AssumePrime = 1;
	end	else if (num==16'd62213) begin
		AssumePrime = 1;
	end	else if (num==16'd62219) begin
		AssumePrime = 1;
	end	else if (num==16'd62233) begin
		AssumePrime = 1;
	end	else if (num==16'd62273) begin
		AssumePrime = 1;
	end	else if (num==16'd62297) begin
		AssumePrime = 1;
	end	else if (num==16'd62299) begin
		AssumePrime = 1;
	end	else if (num==16'd62303) begin
		AssumePrime = 1;
	end	else if (num==16'd62311) begin
		AssumePrime = 1;
	end	else if (num==16'd62323) begin
		AssumePrime = 1;
	end	else if (num==16'd62327) begin
		AssumePrime = 1;
	end	else if (num==16'd62347) begin
		AssumePrime = 1;
	end	else if (num==16'd62351) begin
		AssumePrime = 1;
	end	else if (num==16'd62383) begin
		AssumePrime = 1;
	end	else if (num==16'd62401) begin
		AssumePrime = 1;
	end	else if (num==16'd62417) begin
		AssumePrime = 1;
	end	else if (num==16'd62423) begin
		AssumePrime = 1;
	end	else if (num==16'd62459) begin
		AssumePrime = 1;
	end	else if (num==16'd62467) begin
		AssumePrime = 1;
	end	else if (num==16'd62473) begin
		AssumePrime = 1;
	end	else if (num==16'd62477) begin
		AssumePrime = 1;
	end	else if (num==16'd62483) begin
		AssumePrime = 1;
	end	else if (num==16'd62497) begin
		AssumePrime = 1;
	end	else if (num==16'd62501) begin
		AssumePrime = 1;
	end	else if (num==16'd62507) begin
		AssumePrime = 1;
	end	else if (num==16'd62533) begin
		AssumePrime = 1;
	end	else if (num==16'd62539) begin
		AssumePrime = 1;
	end	else if (num==16'd62549) begin
		AssumePrime = 1;
	end	else if (num==16'd62563) begin
		AssumePrime = 1;
	end	else if (num==16'd62581) begin
		AssumePrime = 1;
	end	else if (num==16'd62591) begin
		AssumePrime = 1;
	end	else if (num==16'd62597) begin
		AssumePrime = 1;
	end	else if (num==16'd62603) begin
		AssumePrime = 1;
	end	else if (num==16'd62617) begin
		AssumePrime = 1;
	end	else if (num==16'd62627) begin
		AssumePrime = 1;
	end	else if (num==16'd62633) begin
		AssumePrime = 1;
	end	else if (num==16'd62639) begin
		AssumePrime = 1;
	end	else if (num==16'd62653) begin
		AssumePrime = 1;
	end	else if (num==16'd62659) begin
		AssumePrime = 1;
	end	else if (num==16'd62683) begin
		AssumePrime = 1;
	end	else if (num==16'd62687) begin
		AssumePrime = 1;
	end	else if (num==16'd62701) begin
		AssumePrime = 1;
	end	else if (num==16'd62723) begin
		AssumePrime = 1;
	end	else if (num==16'd62731) begin
		AssumePrime = 1;
	end	else if (num==16'd62743) begin
		AssumePrime = 1;
	end	else if (num==16'd62753) begin
		AssumePrime = 1;
	end	else if (num==16'd62761) begin
		AssumePrime = 1;
	end	else if (num==16'd62773) begin
		AssumePrime = 1;
	end	else if (num==16'd62791) begin
		AssumePrime = 1;
	end	else if (num==16'd62801) begin
		AssumePrime = 1;
	end	else if (num==16'd62819) begin
		AssumePrime = 1;
	end	else if (num==16'd62827) begin
		AssumePrime = 1;
	end	else if (num==16'd62851) begin
		AssumePrime = 1;
	end	else if (num==16'd62861) begin
		AssumePrime = 1;
	end	else if (num==16'd62869) begin
		AssumePrime = 1;
	end	else if (num==16'd62873) begin
		AssumePrime = 1;
	end	else if (num==16'd62897) begin
		AssumePrime = 1;
	end	else if (num==16'd62903) begin
		AssumePrime = 1;
	end	else if (num==16'd62921) begin
		AssumePrime = 1;
	end	else if (num==16'd62927) begin
		AssumePrime = 1;
	end	else if (num==16'd62929) begin
		AssumePrime = 1;
	end	else if (num==16'd62939) begin
		AssumePrime = 1;
	end	else if (num==16'd62969) begin
		AssumePrime = 1;
	end	else if (num==16'd62971) begin
		AssumePrime = 1;
	end	else if (num==16'd62981) begin
		AssumePrime = 1;
	end	else if (num==16'd62983) begin
		AssumePrime = 1;
	end	else if (num==16'd62987) begin
		AssumePrime = 1;
	end	else if (num==16'd62989) begin
		AssumePrime = 1;
	end	else if (num==16'd63029) begin
		AssumePrime = 1;
	end	else if (num==16'd63031) begin
		AssumePrime = 1;
	end	else if (num==16'd63059) begin
		AssumePrime = 1;
	end	else if (num==16'd63067) begin
		AssumePrime = 1;
	end	else if (num==16'd63073) begin
		AssumePrime = 1;
	end	else if (num==16'd63079) begin
		AssumePrime = 1;
	end	else if (num==16'd63097) begin
		AssumePrime = 1;
	end	else if (num==16'd63103) begin
		AssumePrime = 1;
	end	else if (num==16'd63113) begin
		AssumePrime = 1;
	end	else if (num==16'd63127) begin
		AssumePrime = 1;
	end	else if (num==16'd63131) begin
		AssumePrime = 1;
	end	else if (num==16'd63149) begin
		AssumePrime = 1;
	end	else if (num==16'd63179) begin
		AssumePrime = 1;
	end	else if (num==16'd63197) begin
		AssumePrime = 1;
	end	else if (num==16'd63199) begin
		AssumePrime = 1;
	end	else if (num==16'd63211) begin
		AssumePrime = 1;
	end	else if (num==16'd63241) begin
		AssumePrime = 1;
	end	else if (num==16'd63247) begin
		AssumePrime = 1;
	end	else if (num==16'd63277) begin
		AssumePrime = 1;
	end	else if (num==16'd63281) begin
		AssumePrime = 1;
	end	else if (num==16'd63299) begin
		AssumePrime = 1;
	end	else if (num==16'd63311) begin
		AssumePrime = 1;
	end	else if (num==16'd63313) begin
		AssumePrime = 1;
	end	else if (num==16'd63317) begin
		AssumePrime = 1;
	end	else if (num==16'd63331) begin
		AssumePrime = 1;
	end	else if (num==16'd63337) begin
		AssumePrime = 1;
	end	else if (num==16'd63347) begin
		AssumePrime = 1;
	end	else if (num==16'd63353) begin
		AssumePrime = 1;
	end	else if (num==16'd63361) begin
		AssumePrime = 1;
	end	else if (num==16'd63367) begin
		AssumePrime = 1;
	end	else if (num==16'd63377) begin
		AssumePrime = 1;
	end	else if (num==16'd63389) begin
		AssumePrime = 1;
	end	else if (num==16'd63391) begin
		AssumePrime = 1;
	end	else if (num==16'd63397) begin
		AssumePrime = 1;
	end	else if (num==16'd63409) begin
		AssumePrime = 1;
	end	else if (num==16'd63419) begin
		AssumePrime = 1;
	end	else if (num==16'd63421) begin
		AssumePrime = 1;
	end	else if (num==16'd63439) begin
		AssumePrime = 1;
	end	else if (num==16'd63443) begin
		AssumePrime = 1;
	end	else if (num==16'd63463) begin
		AssumePrime = 1;
	end	else if (num==16'd63467) begin
		AssumePrime = 1;
	end	else if (num==16'd63473) begin
		AssumePrime = 1;
	end	else if (num==16'd63487) begin
		AssumePrime = 1;
	end	else if (num==16'd63493) begin
		AssumePrime = 1;
	end	else if (num==16'd63499) begin
		AssumePrime = 1;
	end	else if (num==16'd63521) begin
		AssumePrime = 1;
	end	else if (num==16'd63527) begin
		AssumePrime = 1;
	end	else if (num==16'd63533) begin
		AssumePrime = 1;
	end	else if (num==16'd63541) begin
		AssumePrime = 1;
	end	else if (num==16'd63559) begin
		AssumePrime = 1;
	end	else if (num==16'd63577) begin
		AssumePrime = 1;
	end	else if (num==16'd63587) begin
		AssumePrime = 1;
	end	else if (num==16'd63589) begin
		AssumePrime = 1;
	end	else if (num==16'd63599) begin
		AssumePrime = 1;
	end	else if (num==16'd63601) begin
		AssumePrime = 1;
	end	else if (num==16'd63607) begin
		AssumePrime = 1;
	end	else if (num==16'd63611) begin
		AssumePrime = 1;
	end	else if (num==16'd63617) begin
		AssumePrime = 1;
	end	else if (num==16'd63629) begin
		AssumePrime = 1;
	end	else if (num==16'd63647) begin
		AssumePrime = 1;
	end	else if (num==16'd63649) begin
		AssumePrime = 1;
	end	else if (num==16'd63659) begin
		AssumePrime = 1;
	end	else if (num==16'd63667) begin
		AssumePrime = 1;
	end	else if (num==16'd63671) begin
		AssumePrime = 1;
	end	else if (num==16'd63689) begin
		AssumePrime = 1;
	end	else if (num==16'd63691) begin
		AssumePrime = 1;
	end	else if (num==16'd63697) begin
		AssumePrime = 1;
	end	else if (num==16'd63703) begin
		AssumePrime = 1;
	end	else if (num==16'd63709) begin
		AssumePrime = 1;
	end	else if (num==16'd63719) begin
		AssumePrime = 1;
	end	else if (num==16'd63727) begin
		AssumePrime = 1;
	end	else if (num==16'd63737) begin
		AssumePrime = 1;
	end	else if (num==16'd63743) begin
		AssumePrime = 1;
	end	else if (num==16'd63761) begin
		AssumePrime = 1;
	end	else if (num==16'd63773) begin
		AssumePrime = 1;
	end	else if (num==16'd63781) begin
		AssumePrime = 1;
	end	else if (num==16'd63793) begin
		AssumePrime = 1;
	end	else if (num==16'd63799) begin
		AssumePrime = 1;
	end	else if (num==16'd63803) begin
		AssumePrime = 1;
	end	else if (num==16'd63809) begin
		AssumePrime = 1;
	end	else if (num==16'd63823) begin
		AssumePrime = 1;
	end	else if (num==16'd63839) begin
		AssumePrime = 1;
	end	else if (num==16'd63841) begin
		AssumePrime = 1;
	end	else if (num==16'd63853) begin
		AssumePrime = 1;
	end	else if (num==16'd63857) begin
		AssumePrime = 1;
	end	else if (num==16'd63863) begin
		AssumePrime = 1;
	end	else if (num==16'd63901) begin
		AssumePrime = 1;
	end	else if (num==16'd63907) begin
		AssumePrime = 1;
	end	else if (num==16'd63913) begin
		AssumePrime = 1;
	end	else if (num==16'd63929) begin
		AssumePrime = 1;
	end	else if (num==16'd63949) begin
		AssumePrime = 1;
	end	else if (num==16'd63977) begin
		AssumePrime = 1;
	end	else if (num==16'd63997) begin
		AssumePrime = 1;
	end	else if (num==16'd64007) begin
		AssumePrime = 1;
	end	else if (num==16'd64013) begin
		AssumePrime = 1;
	end	else if (num==16'd64019) begin
		AssumePrime = 1;
	end	else if (num==16'd64033) begin
		AssumePrime = 1;
	end	else if (num==16'd64037) begin
		AssumePrime = 1;
	end	else if (num==16'd64063) begin
		AssumePrime = 1;
	end	else if (num==16'd64067) begin
		AssumePrime = 1;
	end	else if (num==16'd64081) begin
		AssumePrime = 1;
	end	else if (num==16'd64091) begin
		AssumePrime = 1;
	end	else if (num==16'd64109) begin
		AssumePrime = 1;
	end	else if (num==16'd64123) begin
		AssumePrime = 1;
	end	else if (num==16'd64151) begin
		AssumePrime = 1;
	end	else if (num==16'd64153) begin
		AssumePrime = 1;
	end	else if (num==16'd64157) begin
		AssumePrime = 1;
	end	else if (num==16'd64171) begin
		AssumePrime = 1;
	end	else if (num==16'd64187) begin
		AssumePrime = 1;
	end	else if (num==16'd64189) begin
		AssumePrime = 1;
	end	else if (num==16'd64217) begin
		AssumePrime = 1;
	end	else if (num==16'd64223) begin
		AssumePrime = 1;
	end	else if (num==16'd64231) begin
		AssumePrime = 1;
	end	else if (num==16'd64237) begin
		AssumePrime = 1;
	end	else if (num==16'd64271) begin
		AssumePrime = 1;
	end	else if (num==16'd64279) begin
		AssumePrime = 1;
	end	else if (num==16'd64283) begin
		AssumePrime = 1;
	end	else if (num==16'd64301) begin
		AssumePrime = 1;
	end	else if (num==16'd64303) begin
		AssumePrime = 1;
	end	else if (num==16'd64319) begin
		AssumePrime = 1;
	end	else if (num==16'd64327) begin
		AssumePrime = 1;
	end	else if (num==16'd64333) begin
		AssumePrime = 1;
	end	else if (num==16'd64373) begin
		AssumePrime = 1;
	end	else if (num==16'd64381) begin
		AssumePrime = 1;
	end	else if (num==16'd64399) begin
		AssumePrime = 1;
	end	else if (num==16'd64403) begin
		AssumePrime = 1;
	end	else if (num==16'd64433) begin
		AssumePrime = 1;
	end	else if (num==16'd64439) begin
		AssumePrime = 1;
	end	else if (num==16'd64451) begin
		AssumePrime = 1;
	end	else if (num==16'd64453) begin
		AssumePrime = 1;
	end	else if (num==16'd64483) begin
		AssumePrime = 1;
	end	else if (num==16'd64489) begin
		AssumePrime = 1;
	end	else if (num==16'd64499) begin
		AssumePrime = 1;
	end	else if (num==16'd64513) begin
		AssumePrime = 1;
	end	else if (num==16'd64553) begin
		AssumePrime = 1;
	end	else if (num==16'd64567) begin
		AssumePrime = 1;
	end	else if (num==16'd64577) begin
		AssumePrime = 1;
	end	else if (num==16'd64579) begin
		AssumePrime = 1;
	end	else if (num==16'd64591) begin
		AssumePrime = 1;
	end	else if (num==16'd64601) begin
		AssumePrime = 1;
	end	else if (num==16'd64609) begin
		AssumePrime = 1;
	end	else if (num==16'd64613) begin
		AssumePrime = 1;
	end	else if (num==16'd64621) begin
		AssumePrime = 1;
	end	else if (num==16'd64627) begin
		AssumePrime = 1;
	end	else if (num==16'd64633) begin
		AssumePrime = 1;
	end	else if (num==16'd64661) begin
		AssumePrime = 1;
	end	else if (num==16'd64663) begin
		AssumePrime = 1;
	end	else if (num==16'd64667) begin
		AssumePrime = 1;
	end	else if (num==16'd64679) begin
		AssumePrime = 1;
	end	else if (num==16'd64693) begin
		AssumePrime = 1;
	end	else if (num==16'd64709) begin
		AssumePrime = 1;
	end	else if (num==16'd64717) begin
		AssumePrime = 1;
	end	else if (num==16'd64747) begin
		AssumePrime = 1;
	end	else if (num==16'd64763) begin
		AssumePrime = 1;
	end	else if (num==16'd64781) begin
		AssumePrime = 1;
	end	else if (num==16'd64783) begin
		AssumePrime = 1;
	end	else if (num==16'd64793) begin
		AssumePrime = 1;
	end	else if (num==16'd64811) begin
		AssumePrime = 1;
	end	else if (num==16'd64817) begin
		AssumePrime = 1;
	end	else if (num==16'd64849) begin
		AssumePrime = 1;
	end	else if (num==16'd64853) begin
		AssumePrime = 1;
	end	else if (num==16'd64871) begin
		AssumePrime = 1;
	end	else if (num==16'd64877) begin
		AssumePrime = 1;
	end	else if (num==16'd64879) begin
		AssumePrime = 1;
	end	else if (num==16'd64891) begin
		AssumePrime = 1;
	end	else if (num==16'd64901) begin
		AssumePrime = 1;
	end	else if (num==16'd64919) begin
		AssumePrime = 1;
	end	else if (num==16'd64921) begin
		AssumePrime = 1;
	end	else if (num==16'd64927) begin
		AssumePrime = 1;
	end	else if (num==16'd64937) begin
		AssumePrime = 1;
	end	else if (num==16'd64951) begin
		AssumePrime = 1;
	end	else if (num==16'd64969) begin
		AssumePrime = 1;
	end	else if (num==16'd64997) begin
		AssumePrime = 1;
	end	else if (num==16'd65003) begin
		AssumePrime = 1;
	end	else if (num==16'd65011) begin
		AssumePrime = 1;
	end	else if (num==16'd65027) begin
		AssumePrime = 1;
	end	else if (num==16'd65029) begin
		AssumePrime = 1;
	end	else if (num==16'd65033) begin
		AssumePrime = 1;
	end	else if (num==16'd65053) begin
		AssumePrime = 1;
	end	else if (num==16'd65063) begin
		AssumePrime = 1;
	end	else if (num==16'd65071) begin
		AssumePrime = 1;
	end	else if (num==16'd65089) begin
		AssumePrime = 1;
	end	else if (num==16'd65099) begin
		AssumePrime = 1;
	end	else if (num==16'd65101) begin
		AssumePrime = 1;
	end	else if (num==16'd65111) begin
		AssumePrime = 1;
	end	else if (num==16'd65119) begin
		AssumePrime = 1;
	end	else if (num==16'd65123) begin
		AssumePrime = 1;
	end	else if (num==16'd65129) begin
		AssumePrime = 1;
	end	else if (num==16'd65141) begin
		AssumePrime = 1;
	end	else if (num==16'd65147) begin
		AssumePrime = 1;
	end	else if (num==16'd65167) begin
		AssumePrime = 1;
	end	else if (num==16'd65171) begin
		AssumePrime = 1;
	end	else if (num==16'd65173) begin
		AssumePrime = 1;
	end	else if (num==16'd65179) begin
		AssumePrime = 1;
	end	else if (num==16'd65183) begin
		AssumePrime = 1;
	end	else if (num==16'd65203) begin
		AssumePrime = 1;
	end	else if (num==16'd65213) begin
		AssumePrime = 1;
	end	else if (num==16'd65239) begin
		AssumePrime = 1;
	end	else if (num==16'd65257) begin
		AssumePrime = 1;
	end	else if (num==16'd65267) begin
		AssumePrime = 1;
	end	else if (num==16'd65269) begin
		AssumePrime = 1;
	end	else if (num==16'd65287) begin
		AssumePrime = 1;
	end	else if (num==16'd65293) begin
		AssumePrime = 1;
	end	else if (num==16'd65309) begin
		AssumePrime = 1;
	end	else if (num==16'd65323) begin
		AssumePrime = 1;
	end	else if (num==16'd65327) begin
		AssumePrime = 1;
	end	else if (num==16'd65353) begin
		AssumePrime = 1;
	end	else if (num==16'd65357) begin
		AssumePrime = 1;
	end	else if (num==16'd65371) begin
		AssumePrime = 1;
	end	else if (num==16'd65381) begin
		AssumePrime = 1;
	end	else if (num==16'd65393) begin
		AssumePrime = 1;
	end	else if (num==16'd65407) begin
		AssumePrime = 1;
	end	else if (num==16'd65413) begin
		AssumePrime = 1;
	end	else if (num==16'd65419) begin
		AssumePrime = 1;
	end	else if (num==16'd65423) begin
		AssumePrime = 1;
	end	else if (num==16'd65437) begin
		AssumePrime = 1;
	end	else if (num==16'd65447) begin
		AssumePrime = 1;
	end	else if (num==16'd65449) begin
		AssumePrime = 1;
	end	else if (num==16'd65479) begin
		AssumePrime = 1;
	end	else if (num==16'd65497) begin
		AssumePrime = 1;
	end	else if (num==16'd65519) begin
		AssumePrime = 1;
	end	else if (num==16'd65521) begin
		AssumePrime = 1;
	end
end


endmodule